** sch_path: /home/leo/Projects/IPs/sky130_leo_ip__comparator/xschem/sky130_leo_ip__comparator.sch
.subckt sky130_leo_ip__comparator vdd in_p out_p in_n vss clk_n out_n
*.PININFO out_n:O in_p:I in_n:I vdd:B vss:B clk_n:I out_p:O
XR1 vss net2 vss sky130_fd_pr__res_xhigh_po_2p85 L=25 mult=1 m=1
XM7 comp_p comp_n vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM1 net2 net2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=5 W=1 nf=1 m=1
XM6 comp_n comp_p vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM2 net1 net2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=5 W=10 nf=1 m=1
XM4 comp_p in_n net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=1 m=1
XM3 comp_n in_p net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=1 m=1
XM5 comp_n clk_n comp_p vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
x1 SR_set net4 VSS VSS VDD VDD net3 sky130_fd_sc_hvl__nand2_1
x2 net3 SR_reset VSS VSS VDD VDD net4 sky130_fd_sc_hvl__nand2_1
XM8 SR_reset comp_p vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM9 SR_reset comp_p vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM10 SR_set comp_n vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM11 SR_set comp_n vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
x3 net3 VSS VSS VDD VDD out_p sky130_fd_sc_hvl__buf_4
x4 net4 VSS VSS VDD VDD out_n sky130_fd_sc_hvl__buf_4
.ends
.end
