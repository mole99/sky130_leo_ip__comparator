* NGSPICE file created from sky130_leo_ip__comparator.ext - technology: sky130A

.subckt sky130_leo_ip__comparator VDD IN_P OUT_P IN_N VSS CLK OUT_N
X0 VSS.t15 a_6094_6197# OUT_P.t6 VSS.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1 a_6602_5707# sky130_fd_sc_hvl__buf_4$VAR1_0.A VSS.t36 VSS.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.07875 pd=0.96 as=0.21375 ps=2.07 w=0.75 l=0.5
X2 VDD.t16 a_84_7283.t3 a_1077_8251.t1 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=3 pd=20.6 as=3 ps=20.6 w=10 l=5
X3 sky130_fd_sc_hvl__buf_4$VAR1_0.A sky130_fd_sc_hvl__nand2_1_0.A a_6602_5227# VSS.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.07875 ps=0.96 w=0.75 l=0.5
X4 sky130_fd_sc_hvl__buf_4$VAR1_0.A SR_set VDD.t20 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X5 OUT_P.t1 a_6094_6197# VDD.t12 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VDD.t10 a_6094_6197# OUT_P.t5 VDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 sky130_fd_sc_hvl__nand2_1_0.A SR_reset a_6602_5707# VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.07875 ps=0.96 w=0.75 l=0.5
X8 sky130_fd_sc_hvl__nand2_1_0.A sky130_fd_sc_hvl__buf_4$VAR1_0.A VDD.t37 VDD.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X9 OUT_N.t3 a_6094_4183# VSS.t27 VSS.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 VDD.t3 COMP_N.t3 SR_set VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=10.6 as=1.5 ps=10.6 w=5 l=0.5
X11 VDD.t18 a_1546_691.t3 SR_reset VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=10.6 as=1.5 ps=10.6 w=5 l=0.5
X12 OUT_N.t7 a_6094_4183# VDD.t29 VDD.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 a_6094_4183# sky130_fd_sc_hvl__buf_4$VAR1_0.A VSS.t34 VSS.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X14 VSS.t13 a_6094_6197# OUT_P.t4 VSS.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X15 VSS.t25 a_6094_4183# OUT_N.t2 VSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X16 a_1546_691.t0 COMP_N.t4 VSS.t3 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=1.5 pd=10.6 as=1.5 ps=10.6 w=5 l=0.5
X17 VSS.t31 sky130_fd_sc_hvl__nand2_1_0.A a_6094_6197# VSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X18 a_84_7283.t2 VSS.t29 VSS.t28 sky130_fd_pr__res_xhigh_po_2p85 l=25.12
X19 COMP_N.t1 IN_P.t0 a_1077_8251.t0 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=6 pd=40.6 as=6 ps=40.6 w=20 l=0.5
X20 VDD.t33 sky130_fd_sc_hvl__nand2_1_0.A sky130_fd_sc_hvl__buf_4$VAR1_0.A VDD.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X21 a_6094_4183# sky130_fd_sc_hvl__buf_4$VAR1_0.A VDD.t35 VDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X22 COMP_N.t0 CLK.t0 a_1546_691.t1 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=3 pd=20.6 as=3 ps=20.6 w=10 l=0.5
X23 VDD.t8 a_6094_6197# OUT_P.t2 VDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X24 VDD.t27 a_6094_4183# OUT_N.t6 VDD.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X25 VDD.t1 SR_reset sky130_fd_sc_hvl__nand2_1_0.A VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X26 a_1077_8251.t2 IN_N.t0 a_1546_691.t2 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=6 pd=40.6 as=6 ps=40.6 w=20 l=0.5
X27 SR_reset a_1546_691.t4 VSS.t17 VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X28 VDD.t31 sky130_fd_sc_hvl__nand2_1_0.A a_6094_6197# VDD.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X29 VSS.t23 a_6094_4183# OUT_N.t1 VSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X30 OUT_P.t7 a_6094_6197# VSS.t11 VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X31 OUT_N.t0 a_6094_4183# VSS.t21 VSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X32 VDD.t25 a_6094_4183# OUT_N.t5 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X33 OUT_P.t3 a_6094_6197# VDD.t6 VDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X34 SR_set COMP_N.t5 VSS.t5 VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X35 VDD.t14 a_84_7283.t0 a_84_7283.t1 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=5
X36 OUT_P.t0 a_6094_6197# VSS.t9 VSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X37 a_6602_5227# SR_set VSS.t19 VSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.07875 pd=0.96 as=0.21375 ps=2.07 w=0.75 l=0.5
X38 OUT_N.t4 a_6094_4183# VDD.t23 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X39 VSS.t7 a_1546_691.t5 COMP_N.t2 VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=1.5 pd=10.6 as=1.5 ps=10.6 w=5 l=0.5
R0 OUT_P.n3 OUT_P.n1 272.034
R1 OUT_P.n6 OUT_P.n4 203.779
R2 OUT_P.n3 OUT_P.n2 181.864
R3 OUT_P.n6 OUT_P.n5 105.144
R4 OUT_P OUT_P.n7 24.3048
R5 OUT_P.n5 OUT_P.t4 21.2805
R6 OUT_P.n5 OUT_P.t0 21.2805
R7 OUT_P.n4 OUT_P.t6 21.2805
R8 OUT_P.n4 OUT_P.t7 21.2805
R9 OUT_P.n2 OUT_P.t2 17.8272
R10 OUT_P.n2 OUT_P.t1 17.8272
R11 OUT_P.n1 OUT_P.t5 17.8272
R12 OUT_P.n1 OUT_P.t3 17.8272
R13 OUT_P.n7 OUT_P.n6 17.529
R14 OUT_P.n7 OUT_P.n3 13.7643
R15 OUT_P OUT_P.n0 8.67196
R16 OUT_P.n0 OUT_P 5.93406
R17 OUT_P.n0 OUT_P 4.27305
R18 VSS.n847 VSS.n184 60168.6
R19 VSS.n759 VSS.n327 30007
R20 VSS.n832 VSS.n831 18043
R21 VSS.n831 VSS.n184 17798.2
R22 VSS.n830 VSS.n829 7706.1
R23 VSS.n829 VSS.n828 7400.63
R24 VSS.n829 VSS.n184 6683.24
R25 VSS.n831 VSS.n830 4658.04
R26 VSS.n849 VSS.n181 1529.65
R27 VSS.n834 VSS.n179 1529.65
R28 VSS.n1065 VSS.n1064 1529.65
R29 VSS.n1139 VSS.n19 1529.65
R30 VSS.n739 VSS.n723 1372.26
R31 VSS.n1095 VSS.n40 722.496
R32 VSS.n596 VSS.n551 665.317
R33 VSS.n594 VSS.n553 665.317
R34 VSS.n603 VSS.n541 665.317
R35 VSS.n633 VSS.n545 665.317
R36 VSS.n722 VSS.n343 665.317
R37 VSS.n708 VSS.n353 665.317
R38 VSS.n432 VSS.n394 665.317
R39 VSS.n387 VSS.n349 665.317
R40 VSS.n638 VSS.n458 652.583
R41 VSS.n533 VSS.n460 652.583
R42 VSS.n645 VSS.n447 652.583
R43 VSS.n703 VSS.n451 652.583
R44 VSS.n749 VSS.n748 652.583
R45 VSS.n732 VSS.n341 652.583
R46 VSS.n741 VSS.n339 652.583
R47 VSS.n757 VSS.n331 652.583
R48 VSS.n305 VSS.n293 652.583
R49 VSS.n316 VSS.n315 652.583
R50 VSS.n326 VSS.n283 652.583
R51 VSS.n308 VSS.n292 652.583
R52 VSS.n302 VSS.n293 585
R53 VSS.n301 VSS.n300 585
R54 VSS.n298 VSS.n294 585
R55 VSS.n296 VSS.n295 585
R56 VSS.n292 VSS.n291 585
R57 VSS.n292 VSS.n188 585
R58 VSS.n309 VSS.n308 585
R59 VSS.n308 VSS.n307 585
R60 VSS.n310 VSS.n290 585
R61 VSS.n306 VSS.n290 585
R62 VSS.n312 VSS.n311 585
R63 VSS.n313 VSS.n312 585
R64 VSS.n285 VSS.n283 585
R65 VSS.n283 VSS.n280 585
R66 VSS.n315 VSS.n287 585
R67 VSS.n315 VSS.n280 585
R68 VSS.n314 VSS.n289 585
R69 VSS.n314 VSS.n313 585
R70 VSS.n303 VSS.n288 585
R71 VSS.n306 VSS.n288 585
R72 VSS.n305 VSS.n304 585
R73 VSS.n307 VSS.n305 585
R74 VSS.n317 VSS.n316 585
R75 VSS.n320 VSS.n319 585
R76 VSS.n322 VSS.n321 585
R77 VSS.n324 VSS.n284 585
R78 VSS.n326 VSS.n325 585
R79 VSS.n327 VSS.n326 585
R80 VSS.n769 VSS.n761 585
R81 VSS.n761 VSS.n760 585
R82 VSS.n771 VSS.n770 585
R83 VSS.n772 VSS.n771 585
R84 VSS.n278 VSS.n277 585
R85 VSS.n773 VSS.n278 585
R86 VSS.n776 VSS.n775 585
R87 VSS.n775 VSS.n774 585
R88 VSS.n777 VSS.n262 585
R89 VSS.n279 VSS.n262 585
R90 VSS.n779 VSS.n778 585
R91 VSS.n780 VSS.n779 585
R92 VSS.n260 VSS.n259 585
R93 VSS.n781 VSS.n260 585
R94 VSS.n784 VSS.n783 585
R95 VSS.n783 VSS.n782 585
R96 VSS.n785 VSS.n247 585
R97 VSS.n261 VSS.n247 585
R98 VSS.n787 VSS.n786 585
R99 VSS.n788 VSS.n787 585
R100 VSS.n245 VSS.n244 585
R101 VSS.n789 VSS.n245 585
R102 VSS.n792 VSS.n791 585
R103 VSS.n791 VSS.n790 585
R104 VSS.n793 VSS.n231 585
R105 VSS.n246 VSS.n231 585
R106 VSS.n795 VSS.n794 585
R107 VSS.n796 VSS.n795 585
R108 VSS.n229 VSS.n228 585
R109 VSS.n797 VSS.n229 585
R110 VSS.n800 VSS.n799 585
R111 VSS.n799 VSS.n798 585
R112 VSS.n801 VSS.n224 585
R113 VSS.n230 VSS.n224 585
R114 VSS.n803 VSS.n802 585
R115 VSS.n804 VSS.n803 585
R116 VSS.n222 VSS.n221 585
R117 VSS.n805 VSS.n222 585
R118 VSS.n808 VSS.n807 585
R119 VSS.n807 VSS.n806 585
R120 VSS.n809 VSS.n210 585
R121 VSS.n223 VSS.n210 585
R122 VSS.n811 VSS.n810 585
R123 VSS.n812 VSS.n811 585
R124 VSS.n208 VSS.n207 585
R125 VSS.n813 VSS.n208 585
R126 VSS.n816 VSS.n815 585
R127 VSS.n815 VSS.n814 585
R128 VSS.n817 VSS.n198 585
R129 VSS.n209 VSS.n198 585
R130 VSS.n819 VSS.n818 585
R131 VSS.n820 VSS.n819 585
R132 VSS.n197 VSS.n196 585
R133 VSS.n821 VSS.n197 585
R134 VSS.n824 VSS.n823 585
R135 VSS.n823 VSS.n822 585
R136 VSS.n825 VSS.n190 585
R137 VSS.n190 VSS.n189 585
R138 VSS.n827 VSS.n826 585
R139 VSS.n828 VSS.n827 585
R140 VSS.n722 VSS.n721 585
R141 VSS.n723 VSS.n722 585
R142 VSS.n720 VSS.n344 585
R143 VSS.n344 VSS.n342 585
R144 VSS.n719 VSS.n718 585
R145 VSS.n718 VSS.n717 585
R146 VSS.n347 VSS.n346 585
R147 VSS.n716 VSS.n347 585
R148 VSS.n366 VSS.n365 585
R149 VSS.n365 VSS.n348 585
R150 VSS.n368 VSS.n367 585
R151 VSS.n369 VSS.n368 585
R152 VSS.n364 VSS.n363 585
R153 VSS.n370 VSS.n364 585
R154 VSS.n373 VSS.n372 585
R155 VSS.n372 VSS.n371 585
R156 VSS.n374 VSS.n362 585
R157 VSS.n362 VSS.n361 585
R158 VSS.n376 VSS.n375 585
R159 VSS.n377 VSS.n376 585
R160 VSS.n360 VSS.n359 585
R161 VSS.n378 VSS.n360 585
R162 VSS.n381 VSS.n380 585
R163 VSS.n380 VSS.n379 585
R164 VSS.n382 VSS.n358 585
R165 VSS.n358 VSS.n357 585
R166 VSS.n384 VSS.n383 585
R167 VSS.n385 VSS.n384 585
R168 VSS.n356 VSS.n355 585
R169 VSS.n388 VSS.n387 585
R170 VSS.n750 VSS.n749 585
R171 VSS.n752 VSS.n751 585
R172 VSS.n754 VSS.n753 585
R173 VSS.n755 VSS.n332 585
R174 VSS.n757 VSS.n756 585
R175 VSS.n758 VSS.n757 585
R176 VSS.n333 VSS.n331 585
R177 VSS.n331 VSS.n328 585
R178 VSS.n745 VSS.n744 585
R179 VSS.n746 VSS.n745 585
R180 VSS.n743 VSS.n337 585
R181 VSS.n340 VSS.n337 585
R182 VSS.n742 VSS.n741 585
R183 VSS.n741 VSS.n740 585
R184 VSS.n731 VSS.n341 585
R185 VSS.n740 VSS.n341 585
R186 VSS.n730 VSS.n335 585
R187 VSS.n340 VSS.n335 585
R188 VSS.n747 VSS.n336 585
R189 VSS.n747 VSS.n746 585
R190 VSS.n748 VSS.n334 585
R191 VSS.n748 VSS.n328 585
R192 VSS.n733 VSS.n732 585
R193 VSS.n735 VSS.n726 585
R194 VSS.n737 VSS.n736 585
R195 VSS.n727 VSS.n725 585
R196 VSS.n339 VSS.n338 585
R197 VSS.n739 VSS.n339 585
R198 VSS.n709 VSS.n708 585
R199 VSS.n708 VSS.n707 585
R200 VSS.n710 VSS.n351 585
R201 VSS.n354 VSS.n351 585
R202 VSS.n712 VSS.n711 585
R203 VSS.n713 VSS.n712 585
R204 VSS.n345 VSS.n343 585
R205 VSS.n714 VSS.n343 585
R206 VSS.n432 VSS.n431 585
R207 VSS.n429 VSS.n402 585
R208 VSS.n428 VSS.n427 585
R209 VSS.n426 VSS.n425 585
R210 VSS.n424 VSS.n423 585
R211 VSS.n422 VSS.n421 585
R212 VSS.n420 VSS.n419 585
R213 VSS.n418 VSS.n417 585
R214 VSS.n416 VSS.n415 585
R215 VSS.n414 VSS.n413 585
R216 VSS.n412 VSS.n411 585
R217 VSS.n410 VSS.n409 585
R218 VSS.n408 VSS.n407 585
R219 VSS.n406 VSS.n405 585
R220 VSS.n404 VSS.n403 585
R221 VSS.n353 VSS.n352 585
R222 VSS.n430 VSS.n394 585
R223 VSS.n707 VSS.n394 585
R224 VSS.n393 VSS.n392 585
R225 VSS.n393 VSS.n354 585
R226 VSS.n391 VSS.n350 585
R227 VSS.n713 VSS.n350 585
R228 VSS.n390 VSS.n349 585
R229 VSS.n714 VSS.n349 585
R230 VSS.n597 VSS.n596 585
R231 VSS.n596 VSS.n595 585
R232 VSS.n598 VSS.n549 585
R233 VSS.n552 VSS.n549 585
R234 VSS.n600 VSS.n599 585
R235 VSS.n601 VSS.n600 585
R236 VSS.n546 VSS.n545 585
R237 VSS.n545 VSS.n542 585
R238 VSS.n633 VSS.n632 585
R239 VSS.n631 VSS.n544 585
R240 VSS.n630 VSS.n543 585
R241 VSS.n635 VSS.n543 585
R242 VSS.n629 VSS.n628 585
R243 VSS.n627 VSS.n626 585
R244 VSS.n625 VSS.n624 585
R245 VSS.n623 VSS.n622 585
R246 VSS.n621 VSS.n620 585
R247 VSS.n619 VSS.n618 585
R248 VSS.n617 VSS.n616 585
R249 VSS.n615 VSS.n614 585
R250 VSS.n613 VSS.n612 585
R251 VSS.n611 VSS.n610 585
R252 VSS.n609 VSS.n608 585
R253 VSS.n607 VSS.n606 585
R254 VSS.n605 VSS.n541 585
R255 VSS.n635 VSS.n541 585
R256 VSS.n592 VSS.n553 585
R257 VSS.n591 VSS.n590 585
R258 VSS.n588 VSS.n556 585
R259 VSS.n586 VSS.n585 585
R260 VSS.n584 VSS.n557 585
R261 VSS.n583 VSS.n582 585
R262 VSS.n580 VSS.n558 585
R263 VSS.n578 VSS.n577 585
R264 VSS.n576 VSS.n559 585
R265 VSS.n575 VSS.n574 585
R266 VSS.n572 VSS.n560 585
R267 VSS.n570 VSS.n569 585
R268 VSS.n568 VSS.n561 585
R269 VSS.n567 VSS.n566 585
R270 VSS.n564 VSS.n562 585
R271 VSS.n551 VSS.n550 585
R272 VSS.n594 VSS.n593 585
R273 VSS.n595 VSS.n594 585
R274 VSS.n554 VSS.n547 585
R275 VSS.n552 VSS.n547 585
R276 VSS.n602 VSS.n548 585
R277 VSS.n602 VSS.n601 585
R278 VSS.n604 VSS.n603 585
R279 VSS.n603 VSS.n542 585
R280 VSS.n639 VSS.n638 585
R281 VSS.n638 VSS.n637 585
R282 VSS.n640 VSS.n456 585
R283 VSS.n459 VSS.n456 585
R284 VSS.n642 VSS.n641 585
R285 VSS.n643 VSS.n642 585
R286 VSS.n452 VSS.n451 585
R287 VSS.n451 VSS.n448 585
R288 VSS.n703 VSS.n702 585
R289 VSS.n701 VSS.n450 585
R290 VSS.n700 VSS.n449 585
R291 VSS.n705 VSS.n449 585
R292 VSS.n699 VSS.n698 585
R293 VSS.n697 VSS.n696 585
R294 VSS.n695 VSS.n694 585
R295 VSS.n693 VSS.n692 585
R296 VSS.n691 VSS.n690 585
R297 VSS.n689 VSS.n688 585
R298 VSS.n687 VSS.n686 585
R299 VSS.n685 VSS.n684 585
R300 VSS.n683 VSS.n682 585
R301 VSS.n681 VSS.n680 585
R302 VSS.n679 VSS.n678 585
R303 VSS.n677 VSS.n676 585
R304 VSS.n675 VSS.n674 585
R305 VSS.n673 VSS.n672 585
R306 VSS.n671 VSS.n670 585
R307 VSS.n669 VSS.n668 585
R308 VSS.n667 VSS.n666 585
R309 VSS.n665 VSS.n664 585
R310 VSS.n663 VSS.n662 585
R311 VSS.n661 VSS.n660 585
R312 VSS.n659 VSS.n658 585
R313 VSS.n657 VSS.n656 585
R314 VSS.n655 VSS.n654 585
R315 VSS.n653 VSS.n652 585
R316 VSS.n651 VSS.n650 585
R317 VSS.n649 VSS.n648 585
R318 VSS.n647 VSS.n447 585
R319 VSS.n705 VSS.n447 585
R320 VSS.n533 VSS.n532 585
R321 VSS.n530 VSS.n475 585
R322 VSS.n529 VSS.n528 585
R323 VSS.n527 VSS.n526 585
R324 VSS.n525 VSS.n524 585
R325 VSS.n523 VSS.n522 585
R326 VSS.n521 VSS.n520 585
R327 VSS.n519 VSS.n518 585
R328 VSS.n517 VSS.n516 585
R329 VSS.n515 VSS.n514 585
R330 VSS.n513 VSS.n512 585
R331 VSS.n511 VSS.n510 585
R332 VSS.n509 VSS.n508 585
R333 VSS.n507 VSS.n506 585
R334 VSS.n505 VSS.n504 585
R335 VSS.n503 VSS.n502 585
R336 VSS.n501 VSS.n500 585
R337 VSS.n499 VSS.n498 585
R338 VSS.n497 VSS.n496 585
R339 VSS.n495 VSS.n494 585
R340 VSS.n493 VSS.n492 585
R341 VSS.n491 VSS.n490 585
R342 VSS.n489 VSS.n488 585
R343 VSS.n487 VSS.n486 585
R344 VSS.n485 VSS.n484 585
R345 VSS.n483 VSS.n482 585
R346 VSS.n481 VSS.n480 585
R347 VSS.n479 VSS.n478 585
R348 VSS.n477 VSS.n476 585
R349 VSS.n458 VSS.n457 585
R350 VSS.n531 VSS.n460 585
R351 VSS.n637 VSS.n460 585
R352 VSS.n454 VSS.n453 585
R353 VSS.n459 VSS.n453 585
R354 VSS.n644 VSS.n455 585
R355 VSS.n644 VSS.n643 585
R356 VSS.n646 VSS.n645 585
R357 VSS.n645 VSS.n448 585
R358 VSS.n179 VSS.n178 585
R359 VSS.n180 VSS.n179 585
R360 VSS.n856 VSS.n855 585
R361 VSS.n855 VSS.n854 585
R362 VSS.n857 VSS.n177 585
R363 VSS.n177 VSS.n176 585
R364 VSS.n859 VSS.n858 585
R365 VSS.n860 VSS.n859 585
R366 VSS.n171 VSS.n170 585
R367 VSS.n172 VSS.n171 585
R368 VSS.n868 VSS.n867 585
R369 VSS.n867 VSS.n866 585
R370 VSS.n869 VSS.n169 585
R371 VSS.n169 VSS.n168 585
R372 VSS.n871 VSS.n870 585
R373 VSS.n872 VSS.n871 585
R374 VSS.n163 VSS.n162 585
R375 VSS.n164 VSS.n163 585
R376 VSS.n880 VSS.n879 585
R377 VSS.n879 VSS.n878 585
R378 VSS.n881 VSS.n161 585
R379 VSS.n161 VSS.n160 585
R380 VSS.n883 VSS.n882 585
R381 VSS.n884 VSS.n883 585
R382 VSS.n155 VSS.n154 585
R383 VSS.n156 VSS.n155 585
R384 VSS.n892 VSS.n891 585
R385 VSS.n891 VSS.n890 585
R386 VSS.n893 VSS.n153 585
R387 VSS.n153 VSS.n152 585
R388 VSS.n895 VSS.n894 585
R389 VSS.n896 VSS.n895 585
R390 VSS.n147 VSS.n146 585
R391 VSS.n148 VSS.n147 585
R392 VSS.n904 VSS.n903 585
R393 VSS.n903 VSS.n902 585
R394 VSS.n905 VSS.n145 585
R395 VSS.n145 VSS.n144 585
R396 VSS.n907 VSS.n906 585
R397 VSS.n908 VSS.n907 585
R398 VSS.n139 VSS.n138 585
R399 VSS.n140 VSS.n139 585
R400 VSS.n916 VSS.n915 585
R401 VSS.n915 VSS.n914 585
R402 VSS.n917 VSS.n137 585
R403 VSS.n137 VSS.n136 585
R404 VSS.n919 VSS.n918 585
R405 VSS.n920 VSS.n919 585
R406 VSS.n131 VSS.n130 585
R407 VSS.n132 VSS.n131 585
R408 VSS.n928 VSS.n927 585
R409 VSS.n927 VSS.n926 585
R410 VSS.n929 VSS.n129 585
R411 VSS.n129 VSS.n128 585
R412 VSS.n931 VSS.n930 585
R413 VSS.n932 VSS.n931 585
R414 VSS.n123 VSS.n122 585
R415 VSS.n124 VSS.n123 585
R416 VSS.n940 VSS.n939 585
R417 VSS.n939 VSS.n938 585
R418 VSS.n941 VSS.n121 585
R419 VSS.n121 VSS.n120 585
R420 VSS.n943 VSS.n942 585
R421 VSS.n944 VSS.n943 585
R422 VSS.n115 VSS.n114 585
R423 VSS.n116 VSS.n115 585
R424 VSS.n952 VSS.n951 585
R425 VSS.n951 VSS.n950 585
R426 VSS.n953 VSS.n113 585
R427 VSS.n113 VSS.n112 585
R428 VSS.n955 VSS.n954 585
R429 VSS.n956 VSS.n955 585
R430 VSS.n107 VSS.n106 585
R431 VSS.n108 VSS.n107 585
R432 VSS.n964 VSS.n963 585
R433 VSS.n963 VSS.n962 585
R434 VSS.n965 VSS.n105 585
R435 VSS.n105 VSS.n104 585
R436 VSS.n968 VSS.n967 585
R437 VSS.n969 VSS.n968 585
R438 VSS.n966 VSS.n99 585
R439 VSS.n100 VSS.n99 585
R440 VSS.n976 VSS.n98 585
R441 VSS.n976 VSS.n975 585
R442 VSS.n978 VSS.n977 585
R443 VSS.n977 VSS.n56 585
R444 VSS.n979 VSS.n57 585
R445 VSS.n1054 VSS.n57 585
R446 VSS.n981 VSS.n980 585
R447 VSS.n980 VSS.n58 585
R448 VSS.n982 VSS.n64 585
R449 VSS.n1048 VSS.n64 585
R450 VSS.n983 VSS.n65 585
R451 VSS.n1047 VSS.n65 585
R452 VSS.n984 VSS.n66 585
R453 VSS.n1046 VSS.n66 585
R454 VSS.n986 VSS.n985 585
R455 VSS.n985 VSS.n67 585
R456 VSS.n987 VSS.n71 585
R457 VSS.n1040 VSS.n71 585
R458 VSS.n988 VSS.n72 585
R459 VSS.n1039 VSS.n72 585
R460 VSS.n989 VSS.n73 585
R461 VSS.n1038 VSS.n73 585
R462 VSS.n991 VSS.n990 585
R463 VSS.n990 VSS.n74 585
R464 VSS.n992 VSS.n78 585
R465 VSS.n1032 VSS.n78 585
R466 VSS.n993 VSS.n79 585
R467 VSS.n1031 VSS.n79 585
R468 VSS.n994 VSS.n80 585
R469 VSS.n1030 VSS.n80 585
R470 VSS.n996 VSS.n995 585
R471 VSS.n995 VSS.n81 585
R472 VSS.n997 VSS.n85 585
R473 VSS.n1024 VSS.n85 585
R474 VSS.n998 VSS.n86 585
R475 VSS.n1023 VSS.n86 585
R476 VSS.n999 VSS.n87 585
R477 VSS.n1022 VSS.n87 585
R478 VSS.n1001 VSS.n1000 585
R479 VSS.n1000 VSS.n88 585
R480 VSS.n1002 VSS.n92 585
R481 VSS.n1016 VSS.n92 585
R482 VSS.n1003 VSS.n93 585
R483 VSS.n1015 VSS.n93 585
R484 VSS.n1004 VSS.n94 585
R485 VSS.n1014 VSS.n94 585
R486 VSS.n1005 VSS.n97 585
R487 VSS.n97 VSS.n95 585
R488 VSS.n1007 VSS.n1006 585
R489 VSS.n1008 VSS.n1007 585
R490 VSS.n32 VSS.n31 585
R491 VSS.n33 VSS.n32 585
R492 VSS.n1103 VSS.n1102 585
R493 VSS.n1102 VSS.n1101 585
R494 VSS.n1104 VSS.n30 585
R495 VSS.n34 VSS.n30 585
R496 VSS.n1106 VSS.n1105 585
R497 VSS.n1108 VSS.n29 585
R498 VSS.n1109 VSS.n28 585
R499 VSS.n1109 VSS.n18 585
R500 VSS.n1112 VSS.n1111 585
R501 VSS.n1113 VSS.n27 585
R502 VSS.n1115 VSS.n1114 585
R503 VSS.n1117 VSS.n26 585
R504 VSS.n1120 VSS.n1119 585
R505 VSS.n1121 VSS.n25 585
R506 VSS.n1123 VSS.n1122 585
R507 VSS.n1125 VSS.n24 585
R508 VSS.n1128 VSS.n1127 585
R509 VSS.n1129 VSS.n23 585
R510 VSS.n1131 VSS.n1130 585
R511 VSS.n1133 VSS.n22 585
R512 VSS.n1136 VSS.n1135 585
R513 VSS.n1137 VSS.n19 585
R514 VSS.n850 VSS.n849 585
R515 VSS.n183 VSS.n182 585
R516 VSS.n846 VSS.n845 585
R517 VSS.n847 VSS.n846 585
R518 VSS.n844 VSS.n833 585
R519 VSS.n843 VSS.n842 585
R520 VSS.n841 VSS.n840 585
R521 VSS.n839 VSS.n838 585
R522 VSS.n837 VSS.n836 585
R523 VSS.n835 VSS.n834 585
R524 VSS.n1066 VSS.n1065 585
R525 VSS.n1068 VSS.n1067 585
R526 VSS.n1070 VSS.n1069 585
R527 VSS.n1072 VSS.n1071 585
R528 VSS.n1074 VSS.n1073 585
R529 VSS.n1076 VSS.n1075 585
R530 VSS.n1078 VSS.n1077 585
R531 VSS.n1080 VSS.n1079 585
R532 VSS.n1082 VSS.n1081 585
R533 VSS.n1084 VSS.n1083 585
R534 VSS.n1086 VSS.n1085 585
R535 VSS.n1088 VSS.n1087 585
R536 VSS.n1090 VSS.n1089 585
R537 VSS.n1091 VSS.n49 585
R538 VSS.n1093 VSS.n1092 585
R539 VSS.n39 VSS.n38 585
R540 VSS.n1097 VSS.n1096 585
R541 VSS.n1096 VSS.n1095 585
R542 VSS.n1098 VSS.n36 585
R543 VSS.n36 VSS.n34 585
R544 VSS.n1100 VSS.n1099 585
R545 VSS.n1101 VSS.n1100 585
R546 VSS.n37 VSS.n35 585
R547 VSS.n35 VSS.n33 585
R548 VSS.n1010 VSS.n1009 585
R549 VSS.n1009 VSS.n1008 585
R550 VSS.n1011 VSS.n96 585
R551 VSS.n96 VSS.n95 585
R552 VSS.n1013 VSS.n1012 585
R553 VSS.n1014 VSS.n1013 585
R554 VSS.n91 VSS.n90 585
R555 VSS.n1015 VSS.n91 585
R556 VSS.n1018 VSS.n1017 585
R557 VSS.n1017 VSS.n1016 585
R558 VSS.n1019 VSS.n89 585
R559 VSS.n89 VSS.n88 585
R560 VSS.n1021 VSS.n1020 585
R561 VSS.n1022 VSS.n1021 585
R562 VSS.n84 VSS.n83 585
R563 VSS.n1023 VSS.n84 585
R564 VSS.n1026 VSS.n1025 585
R565 VSS.n1025 VSS.n1024 585
R566 VSS.n1027 VSS.n82 585
R567 VSS.n82 VSS.n81 585
R568 VSS.n1029 VSS.n1028 585
R569 VSS.n1030 VSS.n1029 585
R570 VSS.n77 VSS.n76 585
R571 VSS.n1031 VSS.n77 585
R572 VSS.n1034 VSS.n1033 585
R573 VSS.n1033 VSS.n1032 585
R574 VSS.n1035 VSS.n75 585
R575 VSS.n75 VSS.n74 585
R576 VSS.n1037 VSS.n1036 585
R577 VSS.n1038 VSS.n1037 585
R578 VSS.n70 VSS.n69 585
R579 VSS.n1039 VSS.n70 585
R580 VSS.n1042 VSS.n1041 585
R581 VSS.n1041 VSS.n1040 585
R582 VSS.n1043 VSS.n68 585
R583 VSS.n68 VSS.n67 585
R584 VSS.n1045 VSS.n1044 585
R585 VSS.n1046 VSS.n1045 585
R586 VSS.n63 VSS.n62 585
R587 VSS.n1047 VSS.n63 585
R588 VSS.n1050 VSS.n1049 585
R589 VSS.n1049 VSS.n1048 585
R590 VSS.n1051 VSS.n60 585
R591 VSS.n60 VSS.n58 585
R592 VSS.n1053 VSS.n1052 585
R593 VSS.n1054 VSS.n1053 585
R594 VSS.n61 VSS.n59 585
R595 VSS.n59 VSS.n56 585
R596 VSS.n974 VSS.n973 585
R597 VSS.n975 VSS.n974 585
R598 VSS.n972 VSS.n101 585
R599 VSS.n101 VSS.n100 585
R600 VSS.n971 VSS.n970 585
R601 VSS.n970 VSS.n969 585
R602 VSS.n103 VSS.n102 585
R603 VSS.n104 VSS.n103 585
R604 VSS.n961 VSS.n960 585
R605 VSS.n962 VSS.n961 585
R606 VSS.n959 VSS.n109 585
R607 VSS.n109 VSS.n108 585
R608 VSS.n958 VSS.n957 585
R609 VSS.n957 VSS.n956 585
R610 VSS.n111 VSS.n110 585
R611 VSS.n112 VSS.n111 585
R612 VSS.n949 VSS.n948 585
R613 VSS.n950 VSS.n949 585
R614 VSS.n947 VSS.n117 585
R615 VSS.n117 VSS.n116 585
R616 VSS.n946 VSS.n945 585
R617 VSS.n945 VSS.n944 585
R618 VSS.n119 VSS.n118 585
R619 VSS.n120 VSS.n119 585
R620 VSS.n937 VSS.n936 585
R621 VSS.n938 VSS.n937 585
R622 VSS.n935 VSS.n125 585
R623 VSS.n125 VSS.n124 585
R624 VSS.n934 VSS.n933 585
R625 VSS.n933 VSS.n932 585
R626 VSS.n127 VSS.n126 585
R627 VSS.n128 VSS.n127 585
R628 VSS.n925 VSS.n924 585
R629 VSS.n926 VSS.n925 585
R630 VSS.n923 VSS.n133 585
R631 VSS.n133 VSS.n132 585
R632 VSS.n922 VSS.n921 585
R633 VSS.n921 VSS.n920 585
R634 VSS.n135 VSS.n134 585
R635 VSS.n136 VSS.n135 585
R636 VSS.n913 VSS.n912 585
R637 VSS.n914 VSS.n913 585
R638 VSS.n911 VSS.n141 585
R639 VSS.n141 VSS.n140 585
R640 VSS.n910 VSS.n909 585
R641 VSS.n909 VSS.n908 585
R642 VSS.n143 VSS.n142 585
R643 VSS.n144 VSS.n143 585
R644 VSS.n901 VSS.n900 585
R645 VSS.n902 VSS.n901 585
R646 VSS.n899 VSS.n149 585
R647 VSS.n149 VSS.n148 585
R648 VSS.n898 VSS.n897 585
R649 VSS.n897 VSS.n896 585
R650 VSS.n151 VSS.n150 585
R651 VSS.n152 VSS.n151 585
R652 VSS.n889 VSS.n888 585
R653 VSS.n890 VSS.n889 585
R654 VSS.n887 VSS.n157 585
R655 VSS.n157 VSS.n156 585
R656 VSS.n886 VSS.n885 585
R657 VSS.n885 VSS.n884 585
R658 VSS.n159 VSS.n158 585
R659 VSS.n160 VSS.n159 585
R660 VSS.n877 VSS.n876 585
R661 VSS.n878 VSS.n877 585
R662 VSS.n875 VSS.n165 585
R663 VSS.n165 VSS.n164 585
R664 VSS.n874 VSS.n873 585
R665 VSS.n873 VSS.n872 585
R666 VSS.n167 VSS.n166 585
R667 VSS.n168 VSS.n167 585
R668 VSS.n865 VSS.n864 585
R669 VSS.n866 VSS.n865 585
R670 VSS.n863 VSS.n173 585
R671 VSS.n173 VSS.n172 585
R672 VSS.n862 VSS.n861 585
R673 VSS.n861 VSS.n860 585
R674 VSS.n175 VSS.n174 585
R675 VSS.n176 VSS.n175 585
R676 VSS.n853 VSS.n852 585
R677 VSS.n854 VSS.n853 585
R678 VSS.n851 VSS.n181 585
R679 VSS.n181 VSS.n180 585
R680 VSS.n1139 VSS.n1138 585
R681 VSS.n1140 VSS.n1139 585
R682 VSS.n20 VSS.n16 585
R683 VSS.n1141 VSS.n16 585
R684 VSS.n1144 VSS.n1143 585
R685 VSS.n1143 VSS.n1142 585
R686 VSS.n15 VSS.n13 585
R687 VSS.n17 VSS.n15 585
R688 VSS.n1056 VSS.n1055 585
R689 VSS.n1056 VSS.t28 585
R690 VSS.n1058 VSS.n1057 585
R691 VSS.n1059 VSS.n1058 585
R692 VSS.n53 VSS.n51 585
R693 VSS.n1060 VSS.n51 585
R694 VSS.n1063 VSS.n55 585
R695 VSS.n1063 VSS.n1062 585
R696 VSS.n1064 VSS.n50 585
R697 VSS.n1064 VSS.n41 585
R698 VSS.n830 VSS.n188 558.643
R699 VSS.n760 VSS.n759 550
R700 VSS.n827 VSS.n190 539.294
R701 VSS.n823 VSS.n190 539.294
R702 VSS.n823 VSS.n197 539.294
R703 VSS.n819 VSS.n197 539.294
R704 VSS.n819 VSS.n198 539.294
R705 VSS.n815 VSS.n198 539.294
R706 VSS.n815 VSS.n208 539.294
R707 VSS.n811 VSS.n208 539.294
R708 VSS.n811 VSS.n210 539.294
R709 VSS.n807 VSS.n210 539.294
R710 VSS.n807 VSS.n222 539.294
R711 VSS.n803 VSS.n222 539.294
R712 VSS.n803 VSS.n224 539.294
R713 VSS.n799 VSS.n224 539.294
R714 VSS.n799 VSS.n229 539.294
R715 VSS.n795 VSS.n229 539.294
R716 VSS.n795 VSS.n231 539.294
R717 VSS.n791 VSS.n231 539.294
R718 VSS.n791 VSS.n245 539.294
R719 VSS.n787 VSS.n245 539.294
R720 VSS.n787 VSS.n247 539.294
R721 VSS.n783 VSS.n247 539.294
R722 VSS.n783 VSS.n260 539.294
R723 VSS.n779 VSS.n260 539.294
R724 VSS.n779 VSS.n262 539.294
R725 VSS.n775 VSS.n262 539.294
R726 VSS.n775 VSS.n278 539.294
R727 VSS.n771 VSS.n278 539.294
R728 VSS.n771 VSS.n761 539.294
R729 VSS.n828 VSS.n189 463.159
R730 VSS.n822 VSS.n821 463.159
R731 VSS.n814 VSS.n209 463.159
R732 VSS.n813 VSS.n812 463.159
R733 VSS.n806 VSS.n223 463.159
R734 VSS.n806 VSS.n805 463.159
R735 VSS.n798 VSS.n230 463.159
R736 VSS.n798 VSS.n797 463.159
R737 VSS.n797 VSS.n796 463.159
R738 VSS.n790 VSS.n789 463.159
R739 VSS.n789 VSS.n788 463.159
R740 VSS.n782 VSS.n261 463.159
R741 VSS.n781 VSS.n780 463.159
R742 VSS.n774 VSS.n773 463.159
R743 VSS.n772 VSS.n760 463.159
R744 VSS.n223 VSS.t30 429.387
R745 VSS.n788 VSS.t33 429.387
R746 VSS.t0 VSS.n804 410.089
R747 VSS.n246 VSS.t32 410.089
R748 VSS.n846 VSS.n183 394
R749 VSS.n846 VSS.n833 394
R750 VSS.n842 VSS.n841 394
R751 VSS.n838 VSS.n837 394
R752 VSS.n853 VSS.n181 394
R753 VSS.n853 VSS.n175 394
R754 VSS.n861 VSS.n175 394
R755 VSS.n861 VSS.n173 394
R756 VSS.n865 VSS.n173 394
R757 VSS.n865 VSS.n167 394
R758 VSS.n873 VSS.n167 394
R759 VSS.n873 VSS.n165 394
R760 VSS.n877 VSS.n165 394
R761 VSS.n877 VSS.n159 394
R762 VSS.n885 VSS.n159 394
R763 VSS.n885 VSS.n157 394
R764 VSS.n889 VSS.n157 394
R765 VSS.n889 VSS.n151 394
R766 VSS.n897 VSS.n151 394
R767 VSS.n897 VSS.n149 394
R768 VSS.n901 VSS.n149 394
R769 VSS.n901 VSS.n143 394
R770 VSS.n909 VSS.n143 394
R771 VSS.n909 VSS.n141 394
R772 VSS.n913 VSS.n141 394
R773 VSS.n913 VSS.n135 394
R774 VSS.n921 VSS.n135 394
R775 VSS.n921 VSS.n133 394
R776 VSS.n925 VSS.n133 394
R777 VSS.n925 VSS.n127 394
R778 VSS.n933 VSS.n127 394
R779 VSS.n933 VSS.n125 394
R780 VSS.n937 VSS.n125 394
R781 VSS.n937 VSS.n119 394
R782 VSS.n945 VSS.n119 394
R783 VSS.n945 VSS.n117 394
R784 VSS.n949 VSS.n117 394
R785 VSS.n949 VSS.n111 394
R786 VSS.n957 VSS.n111 394
R787 VSS.n957 VSS.n109 394
R788 VSS.n961 VSS.n109 394
R789 VSS.n961 VSS.n103 394
R790 VSS.n970 VSS.n103 394
R791 VSS.n970 VSS.n101 394
R792 VSS.n974 VSS.n101 394
R793 VSS.n974 VSS.n59 394
R794 VSS.n1053 VSS.n59 394
R795 VSS.n1053 VSS.n60 394
R796 VSS.n1049 VSS.n60 394
R797 VSS.n1049 VSS.n63 394
R798 VSS.n1045 VSS.n63 394
R799 VSS.n1045 VSS.n68 394
R800 VSS.n1041 VSS.n68 394
R801 VSS.n1041 VSS.n70 394
R802 VSS.n1037 VSS.n70 394
R803 VSS.n1037 VSS.n75 394
R804 VSS.n1033 VSS.n75 394
R805 VSS.n1033 VSS.n77 394
R806 VSS.n1029 VSS.n77 394
R807 VSS.n1029 VSS.n82 394
R808 VSS.n1025 VSS.n82 394
R809 VSS.n1025 VSS.n84 394
R810 VSS.n1021 VSS.n84 394
R811 VSS.n1021 VSS.n89 394
R812 VSS.n1017 VSS.n89 394
R813 VSS.n1017 VSS.n91 394
R814 VSS.n1013 VSS.n91 394
R815 VSS.n1013 VSS.n96 394
R816 VSS.n1009 VSS.n96 394
R817 VSS.n1009 VSS.n35 394
R818 VSS.n1100 VSS.n35 394
R819 VSS.n1100 VSS.n36 394
R820 VSS.n1096 VSS.n36 394
R821 VSS.n1096 VSS.n39 394
R822 VSS.n1093 VSS.n49 394
R823 VSS.n1089 VSS.n1088 394
R824 VSS.n1085 VSS.n1084 394
R825 VSS.n1081 VSS.n1080 394
R826 VSS.n1077 VSS.n1076 394
R827 VSS.n1073 VSS.n1072 394
R828 VSS.n1069 VSS.n1068 394
R829 VSS.n1064 VSS.n1063 394
R830 VSS.n1063 VSS.n51 394
R831 VSS.n1058 VSS.n51 394
R832 VSS.n1058 VSS.n1056 394
R833 VSS.n1056 VSS.n15 394
R834 VSS.n1143 VSS.n15 394
R835 VSS.n1143 VSS.n16 394
R836 VSS.n1139 VSS.n16 394
R837 VSS.n855 VSS.n179 394
R838 VSS.n855 VSS.n177 394
R839 VSS.n859 VSS.n177 394
R840 VSS.n859 VSS.n171 394
R841 VSS.n867 VSS.n171 394
R842 VSS.n867 VSS.n169 394
R843 VSS.n871 VSS.n169 394
R844 VSS.n871 VSS.n163 394
R845 VSS.n879 VSS.n163 394
R846 VSS.n879 VSS.n161 394
R847 VSS.n883 VSS.n161 394
R848 VSS.n883 VSS.n155 394
R849 VSS.n891 VSS.n155 394
R850 VSS.n891 VSS.n153 394
R851 VSS.n895 VSS.n153 394
R852 VSS.n895 VSS.n147 394
R853 VSS.n903 VSS.n147 394
R854 VSS.n903 VSS.n145 394
R855 VSS.n907 VSS.n145 394
R856 VSS.n907 VSS.n139 394
R857 VSS.n915 VSS.n139 394
R858 VSS.n915 VSS.n137 394
R859 VSS.n919 VSS.n137 394
R860 VSS.n919 VSS.n131 394
R861 VSS.n927 VSS.n131 394
R862 VSS.n927 VSS.n129 394
R863 VSS.n931 VSS.n129 394
R864 VSS.n931 VSS.n123 394
R865 VSS.n939 VSS.n123 394
R866 VSS.n939 VSS.n121 394
R867 VSS.n943 VSS.n121 394
R868 VSS.n943 VSS.n115 394
R869 VSS.n951 VSS.n115 394
R870 VSS.n951 VSS.n113 394
R871 VSS.n955 VSS.n113 394
R872 VSS.n955 VSS.n107 394
R873 VSS.n963 VSS.n107 394
R874 VSS.n963 VSS.n105 394
R875 VSS.n968 VSS.n105 394
R876 VSS.n968 VSS.n99 394
R877 VSS.n976 VSS.n99 394
R878 VSS.n977 VSS.n976 394
R879 VSS.n977 VSS.n57 394
R880 VSS.n980 VSS.n57 394
R881 VSS.n980 VSS.n64 394
R882 VSS.n65 VSS.n64 394
R883 VSS.n66 VSS.n65 394
R884 VSS.n985 VSS.n66 394
R885 VSS.n985 VSS.n71 394
R886 VSS.n72 VSS.n71 394
R887 VSS.n73 VSS.n72 394
R888 VSS.n990 VSS.n73 394
R889 VSS.n990 VSS.n78 394
R890 VSS.n79 VSS.n78 394
R891 VSS.n80 VSS.n79 394
R892 VSS.n995 VSS.n80 394
R893 VSS.n995 VSS.n85 394
R894 VSS.n86 VSS.n85 394
R895 VSS.n87 VSS.n86 394
R896 VSS.n1000 VSS.n87 394
R897 VSS.n1000 VSS.n92 394
R898 VSS.n93 VSS.n92 394
R899 VSS.n94 VSS.n93 394
R900 VSS.n97 VSS.n94 394
R901 VSS.n1007 VSS.n97 394
R902 VSS.n1007 VSS.n32 394
R903 VSS.n1102 VSS.n32 394
R904 VSS.n1102 VSS.n30 394
R905 VSS.n1106 VSS.n30 394
R906 VSS.n1109 VSS.n1108 394
R907 VSS.n1111 VSS.n1109 394
R908 VSS.n1115 VSS.n27 394
R909 VSS.n1119 VSS.n1117 394
R910 VSS.n1123 VSS.n25 394
R911 VSS.n1127 VSS.n1125 394
R912 VSS.n1131 VSS.n23 394
R913 VSS.n1135 VSS.n1133 394
R914 VSS.n820 VSS.t14 381.14
R915 VSS.n279 VSS.t26 381.14
R916 VSS.t8 VSS.n820 371.491
R917 VSS.t22 VSS.n279 371.491
R918 VSS.n832 VSS.n180 347.438
R919 VSS.n386 VSS.n385 329.171
R920 VSS.n759 VSS.n758 291.808
R921 VSS.n804 VSS.t35 275
R922 VSS.t18 VSS.n246 275
R923 VSS.t12 VSS.n189 265.351
R924 VSS.t20 VSS.n772 265.351
R925 VSS.t10 VSS.n813 255.702
R926 VSS.n782 VSS.t24 255.702
R927 VSS.n299 VSS.n188 244.588
R928 VSS.n297 VSS.n188 244.588
R929 VSS.n327 VSS.n281 244.588
R930 VSS.n327 VSS.n282 244.588
R931 VSS.n758 VSS.n329 244.588
R932 VSS.n758 VSS.n330 244.588
R933 VSS.n739 VSS.n724 244.588
R934 VSS.n739 VSS.n738 244.588
R935 VSS.n706 VSS.n433 244.588
R936 VSS.n706 VSS.n401 244.588
R937 VSS.n706 VSS.n400 244.588
R938 VSS.n706 VSS.n399 244.588
R939 VSS.n706 VSS.n398 244.588
R940 VSS.n706 VSS.n397 244.588
R941 VSS.n706 VSS.n396 244.588
R942 VSS.n706 VSS.n395 244.588
R943 VSS.n635 VSS.n634 244.588
R944 VSS.n635 VSS.n535 244.588
R945 VSS.n635 VSS.n536 244.588
R946 VSS.n635 VSS.n537 244.588
R947 VSS.n635 VSS.n538 244.588
R948 VSS.n635 VSS.n539 244.588
R949 VSS.n635 VSS.n540 244.588
R950 VSS.n589 VSS.n40 244.588
R951 VSS.n587 VSS.n40 244.588
R952 VSS.n581 VSS.n40 244.588
R953 VSS.n579 VSS.n40 244.588
R954 VSS.n573 VSS.n40 244.588
R955 VSS.n571 VSS.n40 244.588
R956 VSS.n565 VSS.n40 244.588
R957 VSS.n563 VSS.n40 244.588
R958 VSS.n705 VSS.n704 244.588
R959 VSS.n705 VSS.n434 244.588
R960 VSS.n705 VSS.n435 244.588
R961 VSS.n705 VSS.n436 244.588
R962 VSS.n705 VSS.n437 244.588
R963 VSS.n705 VSS.n438 244.588
R964 VSS.n705 VSS.n439 244.588
R965 VSS.n705 VSS.n440 244.588
R966 VSS.n705 VSS.n441 244.588
R967 VSS.n705 VSS.n442 244.588
R968 VSS.n705 VSS.n443 244.588
R969 VSS.n705 VSS.n444 244.588
R970 VSS.n705 VSS.n445 244.588
R971 VSS.n705 VSS.n446 244.588
R972 VSS.n636 VSS.n534 244.588
R973 VSS.n636 VSS.n474 244.588
R974 VSS.n636 VSS.n473 244.588
R975 VSS.n636 VSS.n472 244.588
R976 VSS.n636 VSS.n471 244.588
R977 VSS.n636 VSS.n470 244.588
R978 VSS.n636 VSS.n469 244.588
R979 VSS.n636 VSS.n468 244.588
R980 VSS.n636 VSS.n467 244.588
R981 VSS.n636 VSS.n466 244.588
R982 VSS.n636 VSS.n465 244.588
R983 VSS.n636 VSS.n464 244.588
R984 VSS.n636 VSS.n463 244.588
R985 VSS.n636 VSS.n462 244.588
R986 VSS.n636 VSS.n461 244.588
R987 VSS.n478 VSS.n477 229.201
R988 VSS.n482 VSS.n481 229.201
R989 VSS.n486 VSS.n485 229.201
R990 VSS.n490 VSS.n489 229.201
R991 VSS.n494 VSS.n493 229.201
R992 VSS.n498 VSS.n497 229.201
R993 VSS.n502 VSS.n501 229.201
R994 VSS.n506 VSS.n505 229.201
R995 VSS.n510 VSS.n509 229.201
R996 VSS.n514 VSS.n513 229.201
R997 VSS.n518 VSS.n517 229.201
R998 VSS.n522 VSS.n521 229.201
R999 VSS.n526 VSS.n525 229.201
R1000 VSS.n528 VSS.n475 229.201
R1001 VSS.n645 VSS.n644 229.201
R1002 VSS.n644 VSS.n453 229.201
R1003 VSS.n460 VSS.n453 229.201
R1004 VSS.n450 VSS.n449 229.201
R1005 VSS.n698 VSS.n449 229.201
R1006 VSS.n696 VSS.n695 229.201
R1007 VSS.n692 VSS.n691 229.201
R1008 VSS.n688 VSS.n687 229.201
R1009 VSS.n684 VSS.n683 229.201
R1010 VSS.n680 VSS.n679 229.201
R1011 VSS.n676 VSS.n675 229.201
R1012 VSS.n672 VSS.n671 229.201
R1013 VSS.n668 VSS.n667 229.201
R1014 VSS.n664 VSS.n663 229.201
R1015 VSS.n660 VSS.n659 229.201
R1016 VSS.n656 VSS.n655 229.201
R1017 VSS.n652 VSS.n651 229.201
R1018 VSS.n648 VSS.n447 229.201
R1019 VSS.n642 VSS.n451 229.201
R1020 VSS.n642 VSS.n456 229.201
R1021 VSS.n638 VSS.n456 229.201
R1022 VSS.n566 VSS.n564 229.201
R1023 VSS.n570 VSS.n561 229.201
R1024 VSS.n574 VSS.n572 229.201
R1025 VSS.n578 VSS.n559 229.201
R1026 VSS.n582 VSS.n580 229.201
R1027 VSS.n586 VSS.n557 229.201
R1028 VSS.n590 VSS.n588 229.201
R1029 VSS.n603 VSS.n602 229.201
R1030 VSS.n602 VSS.n547 229.201
R1031 VSS.n594 VSS.n547 229.201
R1032 VSS.n544 VSS.n543 229.201
R1033 VSS.n628 VSS.n543 229.201
R1034 VSS.n626 VSS.n625 229.201
R1035 VSS.n622 VSS.n621 229.201
R1036 VSS.n618 VSS.n617 229.201
R1037 VSS.n614 VSS.n613 229.201
R1038 VSS.n610 VSS.n609 229.201
R1039 VSS.n606 VSS.n541 229.201
R1040 VSS.n600 VSS.n545 229.201
R1041 VSS.n600 VSS.n549 229.201
R1042 VSS.n596 VSS.n549 229.201
R1043 VSS.n748 VSS.n747 229.201
R1044 VSS.n747 VSS.n335 229.201
R1045 VSS.n341 VSS.n335 229.201
R1046 VSS.n725 VSS.n339 229.201
R1047 VSS.n737 VSS.n726 229.201
R1048 VSS.n745 VSS.n331 229.201
R1049 VSS.n745 VSS.n337 229.201
R1050 VSS.n741 VSS.n337 229.201
R1051 VSS.n757 VSS.n332 229.201
R1052 VSS.n753 VSS.n752 229.201
R1053 VSS.n712 VSS.n343 229.201
R1054 VSS.n712 VSS.n351 229.201
R1055 VSS.n708 VSS.n351 229.201
R1056 VSS.n405 VSS.n404 229.201
R1057 VSS.n409 VSS.n408 229.201
R1058 VSS.n413 VSS.n412 229.201
R1059 VSS.n417 VSS.n416 229.201
R1060 VSS.n421 VSS.n420 229.201
R1061 VSS.n425 VSS.n424 229.201
R1062 VSS.n427 VSS.n402 229.201
R1063 VSS.n350 VSS.n349 229.201
R1064 VSS.n393 VSS.n350 229.201
R1065 VSS.n394 VSS.n393 229.201
R1066 VSS.n722 VSS.n344 229.201
R1067 VSS.n718 VSS.n344 229.201
R1068 VSS.n718 VSS.n347 229.201
R1069 VSS.n365 VSS.n347 229.201
R1070 VSS.n368 VSS.n365 229.201
R1071 VSS.n368 VSS.n364 229.201
R1072 VSS.n372 VSS.n364 229.201
R1073 VSS.n372 VSS.n362 229.201
R1074 VSS.n376 VSS.n362 229.201
R1075 VSS.n376 VSS.n360 229.201
R1076 VSS.n380 VSS.n360 229.201
R1077 VSS.n380 VSS.n358 229.201
R1078 VSS.n384 VSS.n358 229.201
R1079 VSS.n384 VSS.n356 229.201
R1080 VSS.n305 VSS.n288 229.201
R1081 VSS.n314 VSS.n288 229.201
R1082 VSS.n315 VSS.n314 229.201
R1083 VSS.n326 VSS.n284 229.201
R1084 VSS.n321 VSS.n320 229.201
R1085 VSS.n308 VSS.n290 229.201
R1086 VSS.n312 VSS.n290 229.201
R1087 VSS.n312 VSS.n283 229.201
R1088 VSS.n296 VSS.n292 229.201
R1089 VSS.n300 VSS.n298 229.201
R1090 VSS.n1107 VSS.n18 218.815
R1091 VSS.n1110 VSS.n18 218.815
R1092 VSS.n1116 VSS.n18 218.815
R1093 VSS.n1118 VSS.n18 218.815
R1094 VSS.n1124 VSS.n18 218.815
R1095 VSS.n1126 VSS.n18 218.815
R1096 VSS.n1132 VSS.n18 218.815
R1097 VSS.n1134 VSS.n18 218.815
R1098 VSS.n848 VSS.n847 218.815
R1099 VSS.n847 VSS.n185 218.815
R1100 VSS.n847 VSS.n186 218.815
R1101 VSS.n847 VSS.n187 218.815
R1102 VSS.n1095 VSS.n42 218.815
R1103 VSS.n1095 VSS.n43 218.815
R1104 VSS.n1095 VSS.n44 218.815
R1105 VSS.n1095 VSS.n45 218.815
R1106 VSS.n1095 VSS.n46 218.815
R1107 VSS.n1095 VSS.n47 218.815
R1108 VSS.n1095 VSS.n48 218.815
R1109 VSS.n1095 VSS.n1094 218.815
R1110 VSS.n814 VSS.t10 207.457
R1111 VSS.t24 VSS.n781 207.457
R1112 VSS.n822 VSS.t12 197.808
R1113 VSS.n773 VSS.t20 197.808
R1114 VSS.n230 VSS.t35 188.159
R1115 VSS.n790 VSS.t18 188.159
R1116 VSS.n203 VSS.n202 185
R1117 VSS.n274 VSS.n273 185
R1118 VSS.n1095 VSS.n41 182.07
R1119 VSS.n1140 VSS.n18 182.07
R1120 VSS.n854 VSS.n180 180.351
R1121 VSS.n854 VSS.n176 180.351
R1122 VSS.n860 VSS.n176 180.351
R1123 VSS.n860 VSS.n172 180.351
R1124 VSS.n866 VSS.n172 180.351
R1125 VSS.n866 VSS.n168 180.351
R1126 VSS.n872 VSS.n168 180.351
R1127 VSS.n872 VSS.n164 180.351
R1128 VSS.n878 VSS.n164 180.351
R1129 VSS.n878 VSS.n160 180.351
R1130 VSS.n884 VSS.n160 180.351
R1131 VSS.n884 VSS.n156 180.351
R1132 VSS.n890 VSS.n156 180.351
R1133 VSS.n890 VSS.n152 180.351
R1134 VSS.n896 VSS.n152 180.351
R1135 VSS.n896 VSS.n148 180.351
R1136 VSS.n902 VSS.n148 180.351
R1137 VSS.n902 VSS.n144 180.351
R1138 VSS.n908 VSS.n144 180.351
R1139 VSS.n908 VSS.n140 180.351
R1140 VSS.n914 VSS.n140 180.351
R1141 VSS.n914 VSS.n136 180.351
R1142 VSS.n920 VSS.n136 180.351
R1143 VSS.n920 VSS.n132 180.351
R1144 VSS.n926 VSS.n132 180.351
R1145 VSS.n926 VSS.n128 180.351
R1146 VSS.n932 VSS.n128 180.351
R1147 VSS.n932 VSS.n124 180.351
R1148 VSS.n938 VSS.n124 180.351
R1149 VSS.n938 VSS.n120 180.351
R1150 VSS.n944 VSS.n120 180.351
R1151 VSS.n944 VSS.n116 180.351
R1152 VSS.n950 VSS.n116 180.351
R1153 VSS.n950 VSS.n112 180.351
R1154 VSS.n956 VSS.n112 180.351
R1155 VSS.n956 VSS.n108 180.351
R1156 VSS.n962 VSS.n108 180.351
R1157 VSS.n962 VSS.n104 180.351
R1158 VSS.n969 VSS.n104 180.351
R1159 VSS.n969 VSS.n100 180.351
R1160 VSS.n975 VSS.n100 180.351
R1161 VSS.n975 VSS.n56 180.351
R1162 VSS.n1054 VSS.n58 180.351
R1163 VSS.n1048 VSS.n58 180.351
R1164 VSS.n1048 VSS.n1047 180.351
R1165 VSS.n1047 VSS.n1046 180.351
R1166 VSS.n1046 VSS.n67 180.351
R1167 VSS.n1040 VSS.n67 180.351
R1168 VSS.n1040 VSS.n1039 180.351
R1169 VSS.n1039 VSS.n1038 180.351
R1170 VSS.n1038 VSS.n74 180.351
R1171 VSS.n1032 VSS.n74 180.351
R1172 VSS.n1032 VSS.n1031 180.351
R1173 VSS.n1031 VSS.n1030 180.351
R1174 VSS.n1030 VSS.n81 180.351
R1175 VSS.n1024 VSS.n81 180.351
R1176 VSS.n1024 VSS.n1023 180.351
R1177 VSS.n1023 VSS.n1022 180.351
R1178 VSS.n1022 VSS.n88 180.351
R1179 VSS.n1016 VSS.n88 180.351
R1180 VSS.n1016 VSS.n1015 180.351
R1181 VSS.n1015 VSS.n1014 180.351
R1182 VSS.n1014 VSS.n95 180.351
R1183 VSS.n1008 VSS.n95 180.351
R1184 VSS.n1008 VSS.n33 180.351
R1185 VSS.n1101 VSS.n33 180.351
R1186 VSS.n1101 VSS.n34 180.351
R1187 VSS.n707 VSS.n706 174.845
R1188 VSS.n705 VSS.n448 174.845
R1189 VSS.n637 VSS.n636 174.845
R1190 VSS.n635 VSS.n542 174.845
R1191 VSS.n595 VSS.n40 174.845
R1192 VSS.n706 VSS.n705 173.399
R1193 VSS.n636 VSS.n635 173.399
R1194 VSS.n307 VSS.n188 167.316
R1195 VSS.n327 VSS.n280 167.316
R1196 VSS.n849 VSS.n848 147.374
R1197 VSS.n833 VSS.n185 147.374
R1198 VSS.n841 VSS.n186 147.374
R1199 VSS.n837 VSS.n187 147.374
R1200 VSS.n1094 VSS.n1093 147.374
R1201 VSS.n1089 VSS.n48 147.374
R1202 VSS.n1085 VSS.n47 147.374
R1203 VSS.n1081 VSS.n46 147.374
R1204 VSS.n1077 VSS.n45 147.374
R1205 VSS.n1073 VSS.n44 147.374
R1206 VSS.n1069 VSS.n43 147.374
R1207 VSS.n1065 VSS.n42 147.374
R1208 VSS.n1107 VSS.n1106 147.374
R1209 VSS.n1111 VSS.n1110 147.374
R1210 VSS.n1116 VSS.n1115 147.374
R1211 VSS.n1119 VSS.n1118 147.374
R1212 VSS.n1124 VSS.n1123 147.374
R1213 VSS.n1127 VSS.n1126 147.374
R1214 VSS.n1132 VSS.n1131 147.374
R1215 VSS.n1135 VSS.n1134 147.374
R1216 VSS.n1108 VSS.n1107 147.374
R1217 VSS.n1110 VSS.n27 147.374
R1218 VSS.n1117 VSS.n1116 147.374
R1219 VSS.n1118 VSS.n25 147.374
R1220 VSS.n1125 VSS.n1124 147.374
R1221 VSS.n1126 VSS.n23 147.374
R1222 VSS.n1133 VSS.n1132 147.374
R1223 VSS.n1134 VSS.n19 147.374
R1224 VSS.n848 VSS.n183 147.374
R1225 VSS.n842 VSS.n185 147.374
R1226 VSS.n838 VSS.n186 147.374
R1227 VSS.n834 VSS.n187 147.374
R1228 VSS.n1068 VSS.n42 147.374
R1229 VSS.n1072 VSS.n43 147.374
R1230 VSS.n1076 VSS.n44 147.374
R1231 VSS.n1080 VSS.n45 147.374
R1232 VSS.n1084 VSS.n46 147.374
R1233 VSS.n1088 VSS.n47 147.374
R1234 VSS.n49 VSS.n48 147.374
R1235 VSS.n1094 VSS.n39 147.374
R1236 VSS.n193 VSS.t13 142.501
R1237 VSS.n238 VSS.t36 142.501
R1238 VSS.n254 VSS.t19 142.501
R1239 VSS.n765 VSS.t21 142.501
R1240 VSS.n286 VSS.t17 131.495
R1241 VSS.n729 VSS.t5 131.495
R1242 VSS.n758 VSS.n328 115.388
R1243 VSS.n740 VSS.n739 115.388
R1244 VSS.n714 VSS.n713 104.04
R1245 VSS.n707 VSS.n354 104.04
R1246 VSS.n643 VSS.n448 104.04
R1247 VSS.n637 VSS.n459 104.04
R1248 VSS.n601 VSS.n542 104.04
R1249 VSS.n595 VSS.n552 104.04
R1250 VSS.n387 VSS.n386 102.067
R1251 VSS.n307 VSS.n306 99.5605
R1252 VSS.n313 VSS.n280 99.5605
R1253 VSS.n835 VSS.n178 99.3887
R1254 VSS.n851 VSS.n850 99.3887
R1255 VSS.n1062 VSS.n41 98.2599
R1256 VSS.n1060 VSS.n1059 98.2599
R1257 VSS.n1059 VSS.t28 98.2599
R1258 VSS.t28 VSS.n17 98.2599
R1259 VSS.n1142 VSS.n17 98.2599
R1260 VSS.n1142 VSS.n1141 98.2599
R1261 VSS.n1141 VSS.n1140 98.2599
R1262 VSS.n1138 VSS.n1137 96.3914
R1263 VSS.n477 VSS.n461 95.8286
R1264 VSS.n481 VSS.n462 95.8286
R1265 VSS.n485 VSS.n463 95.8286
R1266 VSS.n489 VSS.n464 95.8286
R1267 VSS.n493 VSS.n465 95.8286
R1268 VSS.n497 VSS.n466 95.8286
R1269 VSS.n501 VSS.n467 95.8286
R1270 VSS.n505 VSS.n468 95.8286
R1271 VSS.n509 VSS.n469 95.8286
R1272 VSS.n513 VSS.n470 95.8286
R1273 VSS.n517 VSS.n471 95.8286
R1274 VSS.n521 VSS.n472 95.8286
R1275 VSS.n525 VSS.n473 95.8286
R1276 VSS.n528 VSS.n474 95.8286
R1277 VSS.n534 VSS.n533 95.8286
R1278 VSS.n704 VSS.n703 95.8286
R1279 VSS.n698 VSS.n434 95.8286
R1280 VSS.n695 VSS.n435 95.8286
R1281 VSS.n691 VSS.n436 95.8286
R1282 VSS.n687 VSS.n437 95.8286
R1283 VSS.n683 VSS.n438 95.8286
R1284 VSS.n679 VSS.n439 95.8286
R1285 VSS.n675 VSS.n440 95.8286
R1286 VSS.n671 VSS.n441 95.8286
R1287 VSS.n667 VSS.n442 95.8286
R1288 VSS.n663 VSS.n443 95.8286
R1289 VSS.n659 VSS.n444 95.8286
R1290 VSS.n655 VSS.n445 95.8286
R1291 VSS.n651 VSS.n446 95.8286
R1292 VSS.n564 VSS.n563 95.8286
R1293 VSS.n565 VSS.n561 95.8286
R1294 VSS.n572 VSS.n571 95.8286
R1295 VSS.n573 VSS.n559 95.8286
R1296 VSS.n580 VSS.n579 95.8286
R1297 VSS.n581 VSS.n557 95.8286
R1298 VSS.n588 VSS.n587 95.8286
R1299 VSS.n589 VSS.n553 95.8286
R1300 VSS.n634 VSS.n633 95.8286
R1301 VSS.n628 VSS.n535 95.8286
R1302 VSS.n625 VSS.n536 95.8286
R1303 VSS.n621 VSS.n537 95.8286
R1304 VSS.n617 VSS.n538 95.8286
R1305 VSS.n613 VSS.n539 95.8286
R1306 VSS.n609 VSS.n540 95.8286
R1307 VSS.n738 VSS.n737 95.8286
R1308 VSS.n732 VSS.n724 95.8286
R1309 VSS.n753 VSS.n330 95.8286
R1310 VSS.n749 VSS.n329 95.8286
R1311 VSS.n404 VSS.n395 95.8286
R1312 VSS.n408 VSS.n396 95.8286
R1313 VSS.n412 VSS.n397 95.8286
R1314 VSS.n416 VSS.n398 95.8286
R1315 VSS.n420 VSS.n399 95.8286
R1316 VSS.n424 VSS.n400 95.8286
R1317 VSS.n427 VSS.n401 95.8286
R1318 VSS.n433 VSS.n432 95.8286
R1319 VSS.n321 VSS.n282 95.8286
R1320 VSS.n316 VSS.n281 95.8286
R1321 VSS.n298 VSS.n297 95.8286
R1322 VSS.n299 VSS.n293 95.8286
R1323 VSS.n300 VSS.n299 95.8286
R1324 VSS.n297 VSS.n296 95.8286
R1325 VSS.n320 VSS.n281 95.8286
R1326 VSS.n284 VSS.n282 95.8286
R1327 VSS.n752 VSS.n329 95.8286
R1328 VSS.n332 VSS.n330 95.8286
R1329 VSS.n726 VSS.n724 95.8286
R1330 VSS.n738 VSS.n725 95.8286
R1331 VSS.n433 VSS.n402 95.8286
R1332 VSS.n425 VSS.n401 95.8286
R1333 VSS.n421 VSS.n400 95.8286
R1334 VSS.n417 VSS.n399 95.8286
R1335 VSS.n413 VSS.n398 95.8286
R1336 VSS.n409 VSS.n397 95.8286
R1337 VSS.n405 VSS.n396 95.8286
R1338 VSS.n395 VSS.n353 95.8286
R1339 VSS.n634 VSS.n544 95.8286
R1340 VSS.n626 VSS.n535 95.8286
R1341 VSS.n622 VSS.n536 95.8286
R1342 VSS.n618 VSS.n537 95.8286
R1343 VSS.n614 VSS.n538 95.8286
R1344 VSS.n610 VSS.n539 95.8286
R1345 VSS.n606 VSS.n540 95.8286
R1346 VSS.n590 VSS.n589 95.8286
R1347 VSS.n587 VSS.n586 95.8286
R1348 VSS.n582 VSS.n581 95.8286
R1349 VSS.n579 VSS.n578 95.8286
R1350 VSS.n574 VSS.n573 95.8286
R1351 VSS.n571 VSS.n570 95.8286
R1352 VSS.n566 VSS.n565 95.8286
R1353 VSS.n563 VSS.n551 95.8286
R1354 VSS.n704 VSS.n450 95.8286
R1355 VSS.n696 VSS.n434 95.8286
R1356 VSS.n692 VSS.n435 95.8286
R1357 VSS.n688 VSS.n436 95.8286
R1358 VSS.n684 VSS.n437 95.8286
R1359 VSS.n680 VSS.n438 95.8286
R1360 VSS.n676 VSS.n439 95.8286
R1361 VSS.n672 VSS.n440 95.8286
R1362 VSS.n668 VSS.n441 95.8286
R1363 VSS.n664 VSS.n442 95.8286
R1364 VSS.n660 VSS.n443 95.8286
R1365 VSS.n656 VSS.n444 95.8286
R1366 VSS.n652 VSS.n445 95.8286
R1367 VSS.n648 VSS.n446 95.8286
R1368 VSS.n534 VSS.n475 95.8286
R1369 VSS.n526 VSS.n474 95.8286
R1370 VSS.n522 VSS.n473 95.8286
R1371 VSS.n518 VSS.n472 95.8286
R1372 VSS.n514 VSS.n471 95.8286
R1373 VSS.n510 VSS.n470 95.8286
R1374 VSS.n506 VSS.n469 95.8286
R1375 VSS.n502 VSS.n468 95.8286
R1376 VSS.n498 VSS.n467 95.8286
R1377 VSS.n494 VSS.n466 95.8286
R1378 VSS.n490 VSS.n465 95.8286
R1379 VSS.n486 VSS.n464 95.8286
R1380 VSS.n482 VSS.n463 95.8286
R1381 VSS.n478 VSS.n462 95.8286
R1382 VSS.n461 VSS.n458 95.8286
R1383 VSS.n1066 VSS.n50 95.0883
R1384 VSS.n216 VSS.n215 92.5005
R1385 VSS.n264 VSS.n263 92.5005
R1386 VSS.n821 VSS.t8 91.6672
R1387 VSS.n774 VSS.t22 91.6672
R1388 VSS.n386 VSS.n356 91.3462
R1389 VSS.t28 VSS.n56 90.1753
R1390 VSS.t28 VSS.n1054 90.1753
R1391 VSS.n209 VSS.t14 82.018
R1392 VSS.n780 VSS.t26 82.018
R1393 VSS.n746 VSS.n328 68.6611
R1394 VSS.n740 VSS.n340 68.6611
R1395 VSS.n723 VSS.n342 68.6611
R1396 VSS.n717 VSS.n342 68.6611
R1397 VSS.n717 VSS.n716 68.6611
R1398 VSS.n369 VSS.n348 68.6611
R1399 VSS.n370 VSS.n369 68.6611
R1400 VSS.n371 VSS.n370 68.6611
R1401 VSS.n371 VSS.n361 68.6611
R1402 VSS.n377 VSS.n361 68.6611
R1403 VSS.n378 VSS.n377 68.6611
R1404 VSS.n379 VSS.n378 68.6611
R1405 VSS.n379 VSS.n357 68.6611
R1406 VSS.n385 VSS.n357 68.6611
R1407 VSS.n847 VSS.n832 63.6533
R1408 VSS.n1061 VSS.n1060 59.2452
R1409 VSS.n805 VSS.t0 53.0707
R1410 VSS.n796 VSS.t32 53.0707
R1411 VSS.n713 VSS.t6 52.0202
R1412 VSS.n354 VSS.t6 52.0202
R1413 VSS.n643 VSS.t1 52.0202
R1414 VSS.n459 VSS.t1 52.0202
R1415 VSS.n601 VSS.t2 52.0202
R1416 VSS.n552 VSS.t2 52.0202
R1417 VSS.n306 VSS.t16 49.7805
R1418 VSS.n313 VSS.t16 49.7805
R1419 VSS.n597 VSS.n550 44.5872
R1420 VSS.n593 VSS.n592 44.5872
R1421 VSS.n605 VSS.n604 44.5872
R1422 VSS.n632 VSS.n546 44.5872
R1423 VSS.n721 VSS.n345 44.5872
R1424 VSS.n709 VSS.n352 44.5872
R1425 VSS.n431 VSS.n430 44.5872
R1426 VSS.n390 VSS.n388 44.5872
R1427 VSS.n639 VSS.n457 43.7338
R1428 VSS.n532 VSS.n531 43.7338
R1429 VSS.n647 VSS.n646 43.7338
R1430 VSS.n702 VSS.n452 43.7338
R1431 VSS.n756 VSS.n333 43.7338
R1432 VSS.n742 VSS.n338 43.7338
R1433 VSS.n750 VSS.n334 43.7338
R1434 VSS.n733 VSS.n731 43.7338
R1435 VSS.n304 VSS.n302 43.7338
R1436 VSS.n317 VSS.n287 43.7338
R1437 VSS.n325 VSS.n285 43.7338
R1438 VSS.n309 VSS.n291 43.7338
R1439 VSS.n715 VSS.n348 42.9134
R1440 VSS.n1062 VSS.n1061 39.0153
R1441 VSS.n826 VSS.n825 36.1417
R1442 VSS.n825 VSS.n824 36.1417
R1443 VSS.n824 VSS.n196 36.1417
R1444 VSS.n818 VSS.n196 36.1417
R1445 VSS.n818 VSS.n817 36.1417
R1446 VSS.n817 VSS.n816 36.1417
R1447 VSS.n816 VSS.n207 36.1417
R1448 VSS.n810 VSS.n207 36.1417
R1449 VSS.n810 VSS.n809 36.1417
R1450 VSS.n809 VSS.n808 36.1417
R1451 VSS.n808 VSS.n221 36.1417
R1452 VSS.n802 VSS.n221 36.1417
R1453 VSS.n802 VSS.n801 36.1417
R1454 VSS.n801 VSS.n800 36.1417
R1455 VSS.n800 VSS.n228 36.1417
R1456 VSS.n794 VSS.n228 36.1417
R1457 VSS.n794 VSS.n793 36.1417
R1458 VSS.n793 VSS.n792 36.1417
R1459 VSS.n792 VSS.n244 36.1417
R1460 VSS.n786 VSS.n244 36.1417
R1461 VSS.n786 VSS.n785 36.1417
R1462 VSS.n785 VSS.n784 36.1417
R1463 VSS.n784 VSS.n259 36.1417
R1464 VSS.n778 VSS.n259 36.1417
R1465 VSS.n778 VSS.n777 36.1417
R1466 VSS.n777 VSS.n776 36.1417
R1467 VSS.n776 VSS.n277 36.1417
R1468 VSS.n770 VSS.n277 36.1417
R1469 VSS.n770 VSS.n769 36.1417
R1470 VSS.n715 VSS.n714 34.6803
R1471 VSS.n746 VSS.t4 34.3308
R1472 VSS.n340 VSS.t4 34.3308
R1473 VSS.n812 VSS.t30 33.7724
R1474 VSS.n261 VSS.t33 33.7724
R1475 VSS.n716 VSS.n715 25.7482
R1476 VSS.n856 VSS.n178 25.6005
R1477 VSS.n857 VSS.n856 25.6005
R1478 VSS.n858 VSS.n857 25.6005
R1479 VSS.n858 VSS.n170 25.6005
R1480 VSS.n868 VSS.n170 25.6005
R1481 VSS.n869 VSS.n868 25.6005
R1482 VSS.n870 VSS.n869 25.6005
R1483 VSS.n870 VSS.n162 25.6005
R1484 VSS.n880 VSS.n162 25.6005
R1485 VSS.n881 VSS.n880 25.6005
R1486 VSS.n882 VSS.n881 25.6005
R1487 VSS.n882 VSS.n154 25.6005
R1488 VSS.n892 VSS.n154 25.6005
R1489 VSS.n893 VSS.n892 25.6005
R1490 VSS.n894 VSS.n893 25.6005
R1491 VSS.n894 VSS.n146 25.6005
R1492 VSS.n904 VSS.n146 25.6005
R1493 VSS.n905 VSS.n904 25.6005
R1494 VSS.n906 VSS.n905 25.6005
R1495 VSS.n906 VSS.n138 25.6005
R1496 VSS.n916 VSS.n138 25.6005
R1497 VSS.n917 VSS.n916 25.6005
R1498 VSS.n918 VSS.n917 25.6005
R1499 VSS.n918 VSS.n130 25.6005
R1500 VSS.n928 VSS.n130 25.6005
R1501 VSS.n929 VSS.n928 25.6005
R1502 VSS.n930 VSS.n929 25.6005
R1503 VSS.n930 VSS.n122 25.6005
R1504 VSS.n940 VSS.n122 25.6005
R1505 VSS.n941 VSS.n940 25.6005
R1506 VSS.n942 VSS.n941 25.6005
R1507 VSS.n942 VSS.n114 25.6005
R1508 VSS.n952 VSS.n114 25.6005
R1509 VSS.n953 VSS.n952 25.6005
R1510 VSS.n954 VSS.n953 25.6005
R1511 VSS.n954 VSS.n106 25.6005
R1512 VSS.n964 VSS.n106 25.6005
R1513 VSS.n965 VSS.n964 25.6005
R1514 VSS.n967 VSS.n965 25.6005
R1515 VSS.n967 VSS.n966 25.6005
R1516 VSS.n966 VSS.n98 25.6005
R1517 VSS.n978 VSS.n98 25.6005
R1518 VSS.n979 VSS.n978 25.6005
R1519 VSS.n981 VSS.n979 25.6005
R1520 VSS.n982 VSS.n981 25.6005
R1521 VSS.n983 VSS.n982 25.6005
R1522 VSS.n984 VSS.n983 25.6005
R1523 VSS.n986 VSS.n984 25.6005
R1524 VSS.n987 VSS.n986 25.6005
R1525 VSS.n988 VSS.n987 25.6005
R1526 VSS.n989 VSS.n988 25.6005
R1527 VSS.n991 VSS.n989 25.6005
R1528 VSS.n992 VSS.n991 25.6005
R1529 VSS.n993 VSS.n992 25.6005
R1530 VSS.n994 VSS.n993 25.6005
R1531 VSS.n996 VSS.n994 25.6005
R1532 VSS.n997 VSS.n996 25.6005
R1533 VSS.n998 VSS.n997 25.6005
R1534 VSS.n999 VSS.n998 25.6005
R1535 VSS.n1001 VSS.n999 25.6005
R1536 VSS.n1002 VSS.n1001 25.6005
R1537 VSS.n1003 VSS.n1002 25.6005
R1538 VSS.n1004 VSS.n1003 25.6005
R1539 VSS.n1005 VSS.n1004 25.6005
R1540 VSS.n1006 VSS.n1005 25.6005
R1541 VSS.n1006 VSS.n31 25.6005
R1542 VSS.n1103 VSS.n31 25.6005
R1543 VSS.n1104 VSS.n1103 25.6005
R1544 VSS.n1105 VSS.n1104 25.6005
R1545 VSS.n1105 VSS.n29 25.6005
R1546 VSS.n29 VSS.n28 25.6005
R1547 VSS.n1112 VSS.n28 25.6005
R1548 VSS.n1113 VSS.n1112 25.6005
R1549 VSS.n1114 VSS.n1113 25.6005
R1550 VSS.n1114 VSS.n26 25.6005
R1551 VSS.n1120 VSS.n26 25.6005
R1552 VSS.n1121 VSS.n1120 25.6005
R1553 VSS.n1122 VSS.n1121 25.6005
R1554 VSS.n1122 VSS.n24 25.6005
R1555 VSS.n1128 VSS.n24 25.6005
R1556 VSS.n1129 VSS.n1128 25.6005
R1557 VSS.n1130 VSS.n1129 25.6005
R1558 VSS.n1130 VSS.n22 25.6005
R1559 VSS.n1136 VSS.n22 25.6005
R1560 VSS.n1137 VSS.n1136 25.6005
R1561 VSS.n850 VSS.n182 25.6005
R1562 VSS.n845 VSS.n182 25.6005
R1563 VSS.n845 VSS.n844 25.6005
R1564 VSS.n844 VSS.n843 25.6005
R1565 VSS.n843 VSS.n840 25.6005
R1566 VSS.n840 VSS.n839 25.6005
R1567 VSS.n839 VSS.n836 25.6005
R1568 VSS.n836 VSS.n835 25.6005
R1569 VSS.n852 VSS.n851 25.6005
R1570 VSS.n852 VSS.n174 25.6005
R1571 VSS.n862 VSS.n174 25.6005
R1572 VSS.n863 VSS.n862 25.6005
R1573 VSS.n864 VSS.n863 25.6005
R1574 VSS.n864 VSS.n166 25.6005
R1575 VSS.n874 VSS.n166 25.6005
R1576 VSS.n875 VSS.n874 25.6005
R1577 VSS.n876 VSS.n875 25.6005
R1578 VSS.n876 VSS.n158 25.6005
R1579 VSS.n886 VSS.n158 25.6005
R1580 VSS.n887 VSS.n886 25.6005
R1581 VSS.n888 VSS.n887 25.6005
R1582 VSS.n888 VSS.n150 25.6005
R1583 VSS.n898 VSS.n150 25.6005
R1584 VSS.n899 VSS.n898 25.6005
R1585 VSS.n900 VSS.n899 25.6005
R1586 VSS.n900 VSS.n142 25.6005
R1587 VSS.n910 VSS.n142 25.6005
R1588 VSS.n911 VSS.n910 25.6005
R1589 VSS.n912 VSS.n911 25.6005
R1590 VSS.n912 VSS.n134 25.6005
R1591 VSS.n922 VSS.n134 25.6005
R1592 VSS.n923 VSS.n922 25.6005
R1593 VSS.n924 VSS.n923 25.6005
R1594 VSS.n924 VSS.n126 25.6005
R1595 VSS.n934 VSS.n126 25.6005
R1596 VSS.n935 VSS.n934 25.6005
R1597 VSS.n936 VSS.n935 25.6005
R1598 VSS.n936 VSS.n118 25.6005
R1599 VSS.n946 VSS.n118 25.6005
R1600 VSS.n947 VSS.n946 25.6005
R1601 VSS.n948 VSS.n947 25.6005
R1602 VSS.n948 VSS.n110 25.6005
R1603 VSS.n958 VSS.n110 25.6005
R1604 VSS.n959 VSS.n958 25.6005
R1605 VSS.n960 VSS.n959 25.6005
R1606 VSS.n960 VSS.n102 25.6005
R1607 VSS.n971 VSS.n102 25.6005
R1608 VSS.n972 VSS.n971 25.6005
R1609 VSS.n973 VSS.n972 25.6005
R1610 VSS.n973 VSS.n61 25.6005
R1611 VSS.n1052 VSS.n61 25.6005
R1612 VSS.n1052 VSS.n1051 25.6005
R1613 VSS.n1051 VSS.n1050 25.6005
R1614 VSS.n1050 VSS.n62 25.6005
R1615 VSS.n1044 VSS.n62 25.6005
R1616 VSS.n1044 VSS.n1043 25.6005
R1617 VSS.n1043 VSS.n1042 25.6005
R1618 VSS.n1042 VSS.n69 25.6005
R1619 VSS.n1036 VSS.n69 25.6005
R1620 VSS.n1036 VSS.n1035 25.6005
R1621 VSS.n1035 VSS.n1034 25.6005
R1622 VSS.n1034 VSS.n76 25.6005
R1623 VSS.n1028 VSS.n76 25.6005
R1624 VSS.n1028 VSS.n1027 25.6005
R1625 VSS.n1027 VSS.n1026 25.6005
R1626 VSS.n1026 VSS.n83 25.6005
R1627 VSS.n1020 VSS.n83 25.6005
R1628 VSS.n1020 VSS.n1019 25.6005
R1629 VSS.n1019 VSS.n1018 25.6005
R1630 VSS.n1018 VSS.n90 25.6005
R1631 VSS.n1012 VSS.n90 25.6005
R1632 VSS.n1012 VSS.n1011 25.6005
R1633 VSS.n1011 VSS.n1010 25.6005
R1634 VSS.n1010 VSS.n37 25.6005
R1635 VSS.n1099 VSS.n37 25.6005
R1636 VSS.n1099 VSS.n1098 25.6005
R1637 VSS.n1098 VSS.n1097 25.6005
R1638 VSS.n1097 VSS.n38 25.6005
R1639 VSS.n1092 VSS.n38 25.6005
R1640 VSS.n1092 VSS.n1091 25.6005
R1641 VSS.n1091 VSS.n1090 25.6005
R1642 VSS.n1090 VSS.n1087 25.6005
R1643 VSS.n1087 VSS.n1086 25.6005
R1644 VSS.n1086 VSS.n1083 25.6005
R1645 VSS.n1083 VSS.n1082 25.6005
R1646 VSS.n1082 VSS.n1079 25.6005
R1647 VSS.n1079 VSS.n1078 25.6005
R1648 VSS.n1078 VSS.n1075 25.6005
R1649 VSS.n1075 VSS.n1074 25.6005
R1650 VSS.n1074 VSS.n1071 25.6005
R1651 VSS.n1071 VSS.n1070 25.6005
R1652 VSS.n1070 VSS.n1067 25.6005
R1653 VSS.n1067 VSS.n1066 25.6005
R1654 VSS.n202 VSS.t9 21.2805
R1655 VSS.n202 VSS.t15 21.2805
R1656 VSS.n215 VSS.t11 21.2805
R1657 VSS.n215 VSS.t31 21.2805
R1658 VSS.n263 VSS.t34 21.2805
R1659 VSS.n263 VSS.t25 21.2805
R1660 VSS.n273 VSS.t27 21.2805
R1661 VSS.n273 VSS.t23 21.2805
R1662 VSS.n1061 VSS.n34 21.2181
R1663 VSS.n389 VSS.t7 18.9504
R1664 VSS.n555 VSS.t3 18.9489
R1665 VSS.n204 VSS.n203 15.5066
R1666 VSS.n274 VSS.n272 15.5066
R1667 VSS.n476 VSS.n457 15.3605
R1668 VSS.n479 VSS.n476 15.3605
R1669 VSS.n480 VSS.n479 15.3605
R1670 VSS.n483 VSS.n480 15.3605
R1671 VSS.n484 VSS.n483 15.3605
R1672 VSS.n487 VSS.n484 15.3605
R1673 VSS.n488 VSS.n487 15.3605
R1674 VSS.n491 VSS.n488 15.3605
R1675 VSS.n492 VSS.n491 15.3605
R1676 VSS.n495 VSS.n492 15.3605
R1677 VSS.n496 VSS.n495 15.3605
R1678 VSS.n499 VSS.n496 15.3605
R1679 VSS.n500 VSS.n499 15.3605
R1680 VSS.n503 VSS.n500 15.3605
R1681 VSS.n504 VSS.n503 15.3605
R1682 VSS.n507 VSS.n504 15.3605
R1683 VSS.n508 VSS.n507 15.3605
R1684 VSS.n511 VSS.n508 15.3605
R1685 VSS.n512 VSS.n511 15.3605
R1686 VSS.n515 VSS.n512 15.3605
R1687 VSS.n516 VSS.n515 15.3605
R1688 VSS.n519 VSS.n516 15.3605
R1689 VSS.n520 VSS.n519 15.3605
R1690 VSS.n523 VSS.n520 15.3605
R1691 VSS.n524 VSS.n523 15.3605
R1692 VSS.n527 VSS.n524 15.3605
R1693 VSS.n529 VSS.n527 15.3605
R1694 VSS.n530 VSS.n529 15.3605
R1695 VSS.n532 VSS.n530 15.3605
R1696 VSS.n455 VSS.n454 15.3605
R1697 VSS.n702 VSS.n701 15.3605
R1698 VSS.n701 VSS.n700 15.3605
R1699 VSS.n700 VSS.n699 15.3605
R1700 VSS.n699 VSS.n697 15.3605
R1701 VSS.n697 VSS.n694 15.3605
R1702 VSS.n694 VSS.n693 15.3605
R1703 VSS.n693 VSS.n690 15.3605
R1704 VSS.n690 VSS.n689 15.3605
R1705 VSS.n689 VSS.n686 15.3605
R1706 VSS.n686 VSS.n685 15.3605
R1707 VSS.n685 VSS.n682 15.3605
R1708 VSS.n682 VSS.n681 15.3605
R1709 VSS.n681 VSS.n678 15.3605
R1710 VSS.n678 VSS.n677 15.3605
R1711 VSS.n677 VSS.n674 15.3605
R1712 VSS.n674 VSS.n673 15.3605
R1713 VSS.n673 VSS.n670 15.3605
R1714 VSS.n670 VSS.n669 15.3605
R1715 VSS.n669 VSS.n666 15.3605
R1716 VSS.n666 VSS.n665 15.3605
R1717 VSS.n665 VSS.n662 15.3605
R1718 VSS.n662 VSS.n661 15.3605
R1719 VSS.n661 VSS.n658 15.3605
R1720 VSS.n658 VSS.n657 15.3605
R1721 VSS.n657 VSS.n654 15.3605
R1722 VSS.n654 VSS.n653 15.3605
R1723 VSS.n653 VSS.n650 15.3605
R1724 VSS.n650 VSS.n649 15.3605
R1725 VSS.n649 VSS.n647 15.3605
R1726 VSS.n641 VSS.n452 15.3605
R1727 VSS.n641 VSS.n640 15.3605
R1728 VSS.n640 VSS.n639 15.3605
R1729 VSS.n562 VSS.n550 15.3605
R1730 VSS.n567 VSS.n562 15.3605
R1731 VSS.n568 VSS.n567 15.3605
R1732 VSS.n569 VSS.n568 15.3605
R1733 VSS.n569 VSS.n560 15.3605
R1734 VSS.n575 VSS.n560 15.3605
R1735 VSS.n576 VSS.n575 15.3605
R1736 VSS.n577 VSS.n576 15.3605
R1737 VSS.n577 VSS.n558 15.3605
R1738 VSS.n583 VSS.n558 15.3605
R1739 VSS.n584 VSS.n583 15.3605
R1740 VSS.n585 VSS.n584 15.3605
R1741 VSS.n585 VSS.n556 15.3605
R1742 VSS.n591 VSS.n556 15.3605
R1743 VSS.n592 VSS.n591 15.3605
R1744 VSS.n554 VSS.n548 15.3605
R1745 VSS.n593 VSS.n554 15.3605
R1746 VSS.n632 VSS.n631 15.3605
R1747 VSS.n631 VSS.n630 15.3605
R1748 VSS.n630 VSS.n629 15.3605
R1749 VSS.n629 VSS.n627 15.3605
R1750 VSS.n627 VSS.n624 15.3605
R1751 VSS.n624 VSS.n623 15.3605
R1752 VSS.n623 VSS.n620 15.3605
R1753 VSS.n620 VSS.n619 15.3605
R1754 VSS.n619 VSS.n616 15.3605
R1755 VSS.n616 VSS.n615 15.3605
R1756 VSS.n615 VSS.n612 15.3605
R1757 VSS.n612 VSS.n611 15.3605
R1758 VSS.n611 VSS.n608 15.3605
R1759 VSS.n608 VSS.n607 15.3605
R1760 VSS.n607 VSS.n605 15.3605
R1761 VSS.n599 VSS.n546 15.3605
R1762 VSS.n599 VSS.n598 15.3605
R1763 VSS.n598 VSS.n597 15.3605
R1764 VSS.n711 VSS.n345 15.3605
R1765 VSS.n711 VSS.n710 15.3605
R1766 VSS.n710 VSS.n709 15.3605
R1767 VSS.n403 VSS.n352 15.3605
R1768 VSS.n406 VSS.n403 15.3605
R1769 VSS.n407 VSS.n406 15.3605
R1770 VSS.n410 VSS.n407 15.3605
R1771 VSS.n411 VSS.n410 15.3605
R1772 VSS.n414 VSS.n411 15.3605
R1773 VSS.n415 VSS.n414 15.3605
R1774 VSS.n418 VSS.n415 15.3605
R1775 VSS.n419 VSS.n418 15.3605
R1776 VSS.n422 VSS.n419 15.3605
R1777 VSS.n423 VSS.n422 15.3605
R1778 VSS.n426 VSS.n423 15.3605
R1779 VSS.n428 VSS.n426 15.3605
R1780 VSS.n429 VSS.n428 15.3605
R1781 VSS.n431 VSS.n429 15.3605
R1782 VSS.n391 VSS.n390 15.3605
R1783 VSS.n392 VSS.n391 15.3605
R1784 VSS.n721 VSS.n720 15.3605
R1785 VSS.n720 VSS.n719 15.3605
R1786 VSS.n719 VSS.n346 15.3605
R1787 VSS.n366 VSS.n346 15.3605
R1788 VSS.n367 VSS.n366 15.3605
R1789 VSS.n367 VSS.n363 15.3605
R1790 VSS.n373 VSS.n363 15.3605
R1791 VSS.n374 VSS.n373 15.3605
R1792 VSS.n375 VSS.n374 15.3605
R1793 VSS.n375 VSS.n359 15.3605
R1794 VSS.n381 VSS.n359 15.3605
R1795 VSS.n382 VSS.n381 15.3605
R1796 VSS.n383 VSS.n382 15.3605
R1797 VSS.n383 VSS.n355 15.3605
R1798 VSS.n388 VSS.n355 15.3605
R1799 VSS.n744 VSS.n333 15.3605
R1800 VSS.n744 VSS.n743 15.3605
R1801 VSS.n743 VSS.n742 15.3605
R1802 VSS.n756 VSS.n755 15.3605
R1803 VSS.n755 VSS.n754 15.3605
R1804 VSS.n754 VSS.n751 15.3605
R1805 VSS.n751 VSS.n750 15.3605
R1806 VSS.n336 VSS.n334 15.3605
R1807 VSS.n730 VSS.n336 15.3605
R1808 VSS.n731 VSS.n730 15.3605
R1809 VSS.n736 VSS.n727 15.3605
R1810 VSS.n736 VSS.n735 15.3605
R1811 VSS.n304 VSS.n303 15.3605
R1812 VSS.n303 VSS.n289 15.3605
R1813 VSS.n289 VSS.n287 15.3605
R1814 VSS.n325 VSS.n324 15.3605
R1815 VSS.n322 VSS.n319 15.3605
R1816 VSS.n310 VSS.n309 15.3605
R1817 VSS.n311 VSS.n310 15.3605
R1818 VSS.n311 VSS.n285 15.3605
R1819 VSS.n295 VSS.n291 15.3605
R1820 VSS.n295 VSS.n294 15.3605
R1821 VSS.n301 VSS.n294 15.3605
R1822 VSS.n302 VSS.n301 15.3605
R1823 VSS.n214 VSS.n213 14.5369
R1824 VSS.n268 VSS.n267 14.5369
R1825 VSS.n766 VSS.n0 14.1005
R1826 VSS.n235 VSS.n233 14.0025
R1827 VSS.n251 VSS.n249 14.0025
R1828 VSS.n217 VSS.n216 13.955
R1829 VSS.n265 VSS.n264 13.955
R1830 VSS.n194 VSS.n193 13.5672
R1831 VSS.n765 VSS.n764 13.5672
R1832 VSS.n239 VSS.n238 13.4801
R1833 VSS.n255 VSS.n254 13.4801
R1834 VSS.n55 VSS.n52 13.0467
R1835 VSS.n54 VSS.n53 12.062
R1836 VSS.n1057 VSS.n11 11.0774
R1837 VSS.n21 VSS.n20 10.5851
R1838 VSS.n1055 VSS.n12 10.0928
R1839 VSS.n1144 VSS.n14 9.6005
R1840 VSS.n21 VSS.n8 9.47358
R1841 VSS.n52 VSS.n9 9.47358
R1842 VSS.n325 VSS.n286 9.40867
R1843 VSS.n826 VSS.n191 9.33401
R1844 VSS.n554 VSS.n7 9.3005
R1845 VSS.n593 VSS.n555 9.3005
R1846 VSS.n391 VSS.n2 9.3005
R1847 VSS.n390 VSS.n389 9.3005
R1848 VSS.n767 VSS.n766 9.3005
R1849 VSS.n267 VSS.n266 9.3005
R1850 VSS.n251 VSS.n250 9.3005
R1851 VSS.n253 VSS.n252 9.3005
R1852 VSS.n235 VSS.n234 9.3005
R1853 VSS.n237 VSS.n236 9.3005
R1854 VSS.n214 VSS.n211 9.3005
R1855 VSS.n769 VSS.n768 9.3005
R1856 VSS.n770 VSS.n762 9.3005
R1857 VSS.n763 VSS.n277 9.3005
R1858 VSS.n776 VSS.n276 9.3005
R1859 VSS.n777 VSS.n271 9.3005
R1860 VSS.n778 VSS.n270 9.3005
R1861 VSS.n269 VSS.n259 9.3005
R1862 VSS.n784 VSS.n258 9.3005
R1863 VSS.n785 VSS.n257 9.3005
R1864 VSS.n786 VSS.n256 9.3005
R1865 VSS.n248 VSS.n244 9.3005
R1866 VSS.n792 VSS.n243 9.3005
R1867 VSS.n793 VSS.n242 9.3005
R1868 VSS.n794 VSS.n241 9.3005
R1869 VSS.n240 VSS.n228 9.3005
R1870 VSS.n800 VSS.n227 9.3005
R1871 VSS.n801 VSS.n226 9.3005
R1872 VSS.n802 VSS.n225 9.3005
R1873 VSS.n232 VSS.n221 9.3005
R1874 VSS.n808 VSS.n220 9.3005
R1875 VSS.n809 VSS.n219 9.3005
R1876 VSS.n810 VSS.n218 9.3005
R1877 VSS.n212 VSS.n207 9.3005
R1878 VSS.n816 VSS.n206 9.3005
R1879 VSS.n817 VSS.n205 9.3005
R1880 VSS.n818 VSS.n199 9.3005
R1881 VSS.n200 VSS.n196 9.3005
R1882 VSS.n824 VSS.n195 9.3005
R1883 VSS.n825 VSS.n192 9.3005
R1884 VSS.n736 VSS.n729 9.3005
R1885 VSS.n54 VSS.n9 9.3005
R1886 VSS.n14 VSS.n8 9.3005
R1887 VSS.n1146 VSS.n11 9.3005
R1888 VSS.n1146 VSS.n12 9.3005
R1889 VSS.n1146 VSS.n10 9.3005
R1890 VSS.n1146 VSS.n1145 9.3005
R1891 VSS.n13 VSS.n10 9.10819
R1892 VSS.n1145 VSS.n13 8.61589
R1893 VSS.n1145 VSS.n1144 8.12358
R1894 VSS.n1055 VSS.n10 7.63127
R1895 VSS.n20 VSS.n14 7.13896
R1896 VSS.n203 VSS.n201 6.6818
R1897 VSS.n275 VSS.n274 6.6818
R1898 VSS.n1057 VSS.n12 6.64665
R1899 VSS.n1138 VSS.n21 6.15435
R1900 VSS.n193 VSS.n191 6.126
R1901 VSS.n53 VSS.n11 5.66204
R1902 VSS.n237 VSS.n235 4.70254
R1903 VSS.n253 VSS.n251 4.70254
R1904 VSS.n55 VSS.n54 4.67742
R1905 VSS.n734 VSS.n733 4.26392
R1906 VSS.n318 VSS.n317 4.26392
R1907 VSS.n728 VSS.n338 4.24278
R1908 VSS.n646 VSS.n4 4.23905
R1909 VSS.n531 VSS.n5 4.23905
R1910 VSS.n604 VSS.n6 4.23905
R1911 VSS.n430 VSS.n3 4.23905
R1912 VSS.n323 VSS.n322 4.20736
R1913 VSS.n324 VSS.n323 4.20736
R1914 VSS.n455 VSS.n4 4.19541
R1915 VSS.n454 VSS.n5 4.19541
R1916 VSS.n548 VSS.n6 4.19541
R1917 VSS.n392 VSS.n3 4.19541
R1918 VSS.n728 VSS.n727 4.194
R1919 VSS.n735 VSS.n734 4.18603
R1920 VSS.n319 VSS.n318 4.18603
R1921 VSS.n286 VSS.n1 3.79088
R1922 VSS VSS.n1151 3.7228
R1923 VSS.n52 VSS.n50 3.69281
R1924 VSS.n318 VSS.n286 2.68062
R1925 VSS.n734 VSS.n729 2.68062
R1926 VSS.n1147 VSS.n6 2.63153
R1927 VSS.n1149 VSS.n3 2.63018
R1928 VSS.n1148 VSS.n4 2.6154
R1929 VSS.n1148 VSS.n5 2.6154
R1930 VSS.n729 VSS.n728 2.56926
R1931 VSS.n323 VSS.n286 2.54782
R1932 VSS.n1151 VSS.n1 1.16176
R1933 VSS.n1147 VSS.n1146 0.715574
R1934 VSS.n216 VSS.n214 0.582318
R1935 VSS.n267 VSS.n264 0.582318
R1936 VSS.n766 VSS.n765 0.533833
R1937 VSS.n238 VSS.n237 0.522949
R1938 VSS.n254 VSS.n253 0.522949
R1939 VSS.n1146 VSS.t29 0.474942
R1940 VSS.n1150 VSS 0.34193
R1941 VSS.n1150 VSS.n1149 0.20975
R1942 VSS.n729 VSS.n1 0.181722
R1943 VSS.n1148 VSS.n1147 0.148
R1944 VSS.n1149 VSS.n1148 0.14775
R1945 VSS.n555 VSS.n7 0.0972742
R1946 VSS.n389 VSS.n2 0.0972742
R1947 VSS.n1151 VSS.n1150 0.091
R1948 VSS.n200 VSS.n195 0.0815811
R1949 VSS.n206 VSS.n205 0.0815811
R1950 VSS.n219 VSS.n218 0.0815811
R1951 VSS.n232 VSS.n220 0.0815811
R1952 VSS.n241 VSS.n240 0.0815811
R1953 VSS.n257 VSS.n256 0.0815811
R1954 VSS.n270 VSS.n269 0.0815811
R1955 VSS.n763 VSS.n276 0.0815811
R1956 VSS.n233 VSS.n232 0.067223
R1957 VSS.n249 VSS.n241 0.067223
R1958 VSS.n217 VSS.n211 0.0613108
R1959 VSS.n266 VSS.n265 0.0613108
R1960 VSS.n204 VSS.n199 0.0553986
R1961 VSS.n236 VSS.n227 0.0553986
R1962 VSS.n252 VSS.n248 0.0553986
R1963 VSS.n272 VSS.n271 0.0553986
R1964 VSS.n768 VSS.n767 0.0553986
R1965 VSS.n201 VSS.n200 0.05397
R1966 VSS.n276 VSS.n275 0.05397
R1967 VSS.n192 VSS.n191 0.0489446
R1968 VSS.n195 VSS.n194 0.0469527
R1969 VSS.n213 VSS.n212 0.0469527
R1970 VSS.n234 VSS.n225 0.0469527
R1971 VSS.n250 VSS.n242 0.0469527
R1972 VSS.n268 VSS.n258 0.0469527
R1973 VSS.n764 VSS.n763 0.0469527
R1974 VSS VSS.n219 0.0410405
R1975 VSS.n220 VSS 0.0410405
R1976 VSS.n240 VSS 0.0410405
R1977 VSS.n256 VSS 0.0410405
R1978 VSS.n194 VSS.n192 0.0351284
R1979 VSS.n213 VSS.n206 0.0351284
R1980 VSS.n234 VSS.n226 0.0351284
R1981 VSS VSS.n239 0.0351284
R1982 VSS.n250 VSS.n243 0.0351284
R1983 VSS VSS.n255 0.0351284
R1984 VSS.n269 VSS.n268 0.0351284
R1985 VSS.n764 VSS.n762 0.0351284
R1986 VSS VSS.n0 0.0351284
R1987 VSS.n1149 VSS.n2 0.0341021
R1988 VSS.n1147 VSS.n7 0.0327581
R1989 VSS.n201 VSS.n199 0.0289669
R1990 VSS.n275 VSS.n271 0.0289669
R1991 VSS.n205 VSS.n204 0.0266824
R1992 VSS.n236 VSS.n226 0.0266824
R1993 VSS.n252 VSS.n243 0.0266824
R1994 VSS.n272 VSS.n270 0.0266824
R1995 VSS.n767 VSS.n762 0.0266824
R1996 VSS.n212 VSS.n211 0.0148581
R1997 VSS.n233 VSS.n225 0.0148581
R1998 VSS.n249 VSS.n242 0.0148581
R1999 VSS.n266 VSS.n258 0.0148581
R2000 VSS.n1146 VSS.n9 0.00771154
R2001 VSS.n218 VSS.n217 0.00641216
R2002 VSS.n239 VSS.n227 0.00641216
R2003 VSS.n255 VSS.n248 0.00641216
R2004 VSS.n265 VSS.n257 0.00641216
R2005 VSS.n768 VSS.n0 0.00641216
R2006 VSS.n1146 VSS.n8 0.00530769
R2007 a_84_7283.n64 a_84_7283.t1 354.592
R2008 a_84_7283.n20 a_84_7283.n19 152
R2009 a_84_7283.n34 a_84_7283.n33 152
R2010 a_84_7283.n35 a_84_7283.n18 152
R2011 a_84_7283.n38 a_84_7283.n37 152
R2012 a_84_7283.n36 a_84_7283.n12 152
R2013 a_84_7283.n48 a_84_7283.n47 152
R2014 a_84_7283.n49 a_84_7283.n10 152
R2015 a_84_7283.n51 a_84_7283.n50 152
R2016 a_84_7283.n4 a_84_7283.n3 152
R2017 a_84_7283.n61 a_84_7283.n60 152
R2018 a_84_7283.n58 a_84_7283.n56 152
R2019 a_84_7283.n55 a_84_7283.n6 152
R2020 a_84_7283.n54 a_84_7283.n53 152
R2021 a_84_7283.n8 a_84_7283.n7 152
R2022 a_84_7283.n45 a_84_7283.n44 152
R2023 a_84_7283.n42 a_84_7283.n14 152
R2024 a_84_7283.n41 a_84_7283.n40 152
R2025 a_84_7283.n16 a_84_7283.n15 152
R2026 a_84_7283.n31 a_84_7283.n30 152
R2027 a_84_7283.n29 a_84_7283.n22 152
R2028 a_84_7283.n24 a_84_7283.n19 109.918
R2029 a_84_7283.n62 a_84_7283.n61 109.918
R2030 a_84_7283.n29 a_84_7283.n28 109.918
R2031 a_84_7283.n56 a_84_7283.n1 109.918
R2032 a_84_7283.n43 a_84_7283.t3 48.2005
R2033 a_84_7283.n34 a_84_7283.n19 32.7401
R2034 a_84_7283.n35 a_84_7283.n34 32.7401
R2035 a_84_7283.n37 a_84_7283.n35 32.7401
R2036 a_84_7283.n37 a_84_7283.n36 32.7401
R2037 a_84_7283.n49 a_84_7283.n48 32.7401
R2038 a_84_7283.n50 a_84_7283.n49 32.7401
R2039 a_84_7283.n50 a_84_7283.n3 32.7401
R2040 a_84_7283.n61 a_84_7283.n3 32.7401
R2041 a_84_7283.n30 a_84_7283.n29 32.7401
R2042 a_84_7283.n30 a_84_7283.n15 32.7401
R2043 a_84_7283.n41 a_84_7283.n15 32.7401
R2044 a_84_7283.n42 a_84_7283.n41 32.7401
R2045 a_84_7283.n44 a_84_7283.n7 32.7401
R2046 a_84_7283.n54 a_84_7283.n7 32.7401
R2047 a_84_7283.n55 a_84_7283.n54 32.7401
R2048 a_84_7283.n56 a_84_7283.n55 32.7401
R2049 a_84_7283.n25 a_84_7283.n20 27.1064
R2050 a_84_7283.n33 a_84_7283.n20 27.1064
R2051 a_84_7283.n33 a_84_7283.n18 27.1064
R2052 a_84_7283.n38 a_84_7283.n18 27.1064
R2053 a_84_7283.n38 a_84_7283.n12 27.1064
R2054 a_84_7283.n47 a_84_7283.n12 27.1064
R2055 a_84_7283.n47 a_84_7283.n10 27.1064
R2056 a_84_7283.n51 a_84_7283.n10 27.1064
R2057 a_84_7283.n51 a_84_7283.n4 27.1064
R2058 a_84_7283.n60 a_84_7283.n4 27.1064
R2059 a_84_7283.n60 a_84_7283.n2 27.1064
R2060 a_84_7283.n27 a_84_7283.n22 27.1064
R2061 a_84_7283.n31 a_84_7283.n22 27.1064
R2062 a_84_7283.n31 a_84_7283.n16 27.1064
R2063 a_84_7283.n40 a_84_7283.n16 27.1064
R2064 a_84_7283.n40 a_84_7283.n14 27.1064
R2065 a_84_7283.n45 a_84_7283.n14 27.1064
R2066 a_84_7283.n45 a_84_7283.n8 27.1064
R2067 a_84_7283.n53 a_84_7283.n8 27.1064
R2068 a_84_7283.n53 a_84_7283.n6 27.1064
R2069 a_84_7283.n58 a_84_7283.n6 27.1064
R2070 a_84_7283.n58 a_84_7283.n57 27.1064
R2071 a_84_7283.n24 a_84_7283.n23 23.0638
R2072 a_84_7283.n63 a_84_7283.n62 23.0638
R2073 a_84_7283.n28 a_84_7283.n23 23.0638
R2074 a_84_7283.n63 a_84_7283.n1 23.0638
R2075 a_84_7283.n36 a_84_7283.n11 16.3703
R2076 a_84_7283.n48 a_84_7283.n11 16.3703
R2077 a_84_7283.n43 a_84_7283.n42 16.3703
R2078 a_84_7283.n44 a_84_7283.n43 16.3703
R2079 a_84_7283.n25 a_84_7283.n24 11.3247
R2080 a_84_7283.n62 a_84_7283.n2 11.3247
R2081 a_84_7283.n57 a_84_7283.n1 11.3247
R2082 a_84_7283.n28 a_84_7283.n27 11.3247
R2083 a_84_7283.n57 a_84_7283.n0 9.3005
R2084 a_84_7283.n59 a_84_7283.n58 9.3005
R2085 a_84_7283.n6 a_84_7283.n5 9.3005
R2086 a_84_7283.n53 a_84_7283.n52 9.3005
R2087 a_84_7283.n9 a_84_7283.n8 9.3005
R2088 a_84_7283.n46 a_84_7283.n45 9.3005
R2089 a_84_7283.n14 a_84_7283.n13 9.3005
R2090 a_84_7283.n40 a_84_7283.n39 9.3005
R2091 a_84_7283.n17 a_84_7283.n16 9.3005
R2092 a_84_7283.n32 a_84_7283.n31 9.3005
R2093 a_84_7283.n22 a_84_7283.n21 9.3005
R2094 a_84_7283.n27 a_84_7283.n26 9.3005
R2095 a_84_7283.n2 a_84_7283.n0 9.3005
R2096 a_84_7283.n60 a_84_7283.n59 9.3005
R2097 a_84_7283.n5 a_84_7283.n4 9.3005
R2098 a_84_7283.n52 a_84_7283.n51 9.3005
R2099 a_84_7283.n10 a_84_7283.n9 9.3005
R2100 a_84_7283.n47 a_84_7283.n46 9.3005
R2101 a_84_7283.n13 a_84_7283.n12 9.3005
R2102 a_84_7283.n39 a_84_7283.n38 9.3005
R2103 a_84_7283.n18 a_84_7283.n17 9.3005
R2104 a_84_7283.n33 a_84_7283.n32 9.3005
R2105 a_84_7283.n21 a_84_7283.n20 9.3005
R2106 a_84_7283.n26 a_84_7283.n25 9.3005
R2107 a_84_7283.n11 a_84_7283.t0 4.8205
R2108 a_84_7283.t2 a_84_7283.n64 0.874408
R2109 a_84_7283.n64 a_84_7283.n63 0.60984
R2110 a_84_7283.n26 a_84_7283.n23 0.0174811
R2111 a_84_7283.n26 a_84_7283.n21 0.0174811
R2112 a_84_7283.n32 a_84_7283.n21 0.0174811
R2113 a_84_7283.n32 a_84_7283.n17 0.0174811
R2114 a_84_7283.n39 a_84_7283.n17 0.0174811
R2115 a_84_7283.n39 a_84_7283.n13 0.0174811
R2116 a_84_7283.n46 a_84_7283.n13 0.0174811
R2117 a_84_7283.n46 a_84_7283.n9 0.0174811
R2118 a_84_7283.n52 a_84_7283.n9 0.0174811
R2119 a_84_7283.n52 a_84_7283.n5 0.0174811
R2120 a_84_7283.n59 a_84_7283.n5 0.0174811
R2121 a_84_7283.n59 a_84_7283.n0 0.0174811
R2122 a_84_7283.n63 a_84_7283.n0 0.0174811
R2123 a_1077_8251.n73 a_1077_8251.n8 53.1865
R2124 a_1077_8251.n73 a_1077_8251.n57 285.877
R2125 a_1077_8251.n73 a_1077_8251.n58 285.877
R2126 a_1077_8251.n73 a_1077_8251.n59 285.877
R2127 a_1077_8251.n73 a_1077_8251.n60 285.877
R2128 a_1077_8251.n73 a_1077_8251.n61 285.877
R2129 a_1077_8251.n73 a_1077_8251.n62 285.877
R2130 a_1077_8251.n73 a_1077_8251.n63 285.877
R2131 a_1077_8251.n73 a_1077_8251.n64 285.877
R2132 a_1077_8251.n73 a_1077_8251.n65 285.877
R2133 a_1077_8251.n73 a_1077_8251.n66 285.877
R2134 a_1077_8251.n73 a_1077_8251.n67 285.877
R2135 a_1077_8251.n73 a_1077_8251.n68 285.877
R2136 a_1077_8251.n73 a_1077_8251.n69 285.877
R2137 a_1077_8251.n73 a_1077_8251.n70 285.877
R2138 a_1077_8251.n73 a_1077_8251.n71 285.877
R2139 a_1077_8251.n73 a_1077_8251.n72 285.877
R2140 a_1077_8251.n36 a_1077_8251.n37 285.877
R2141 a_1077_8251.n36 a_1077_8251.n38 285.877
R2142 a_1077_8251.n36 a_1077_8251.n39 285.877
R2143 a_1077_8251.n36 a_1077_8251.n40 285.877
R2144 a_1077_8251.n36 a_1077_8251.n41 285.877
R2145 a_1077_8251.n36 a_1077_8251.n42 285.877
R2146 a_1077_8251.n36 a_1077_8251.n43 285.877
R2147 a_1077_8251.n36 a_1077_8251.n44 285.877
R2148 a_1077_8251.n36 a_1077_8251.n45 285.877
R2149 a_1077_8251.n36 a_1077_8251.n46 285.877
R2150 a_1077_8251.n36 a_1077_8251.n47 285.877
R2151 a_1077_8251.n36 a_1077_8251.n48 285.877
R2152 a_1077_8251.n36 a_1077_8251.n49 285.877
R2153 a_1077_8251.n36 a_1077_8251.n50 285.877
R2154 a_1077_8251.n36 a_1077_8251.n51 285.877
R2155 a_1077_8251.n36 a_1077_8251.n52 285.877
R2156 a_1077_8251.n36 a_1077_8251.n11 48.7551
R2157 a_1077_8251.n53 a_1077_8251.n8 33.502
R2158 a_1077_8251.n59 a_1077_8251.n13 18.7629
R2159 a_1077_8251.n63 a_1077_8251.n15 18.7629
R2160 a_1077_8251.n55 a_1077_8251.n54 27.1064
R2161 a_1077_8251.n67 a_1077_8251.n17 18.7629
R2162 a_1077_8251.n71 a_1077_8251.n19 18.7629
R2163 a_1077_8251.n10 a_1077_8251.n56 33.5713
R2164 a_1077_8251.n37 a_1077_8251.n34 18.7629
R2165 a_1077_8251.n12 a_1077_8251.n39 18.7629
R2166 a_1077_8251.n39 a_1077_8251.n32 18.7629
R2167 a_1077_8251.n40 a_1077_8251.n6 18.7629
R2168 a_1077_8251.n41 a_1077_8251.n30 18.7629
R2169 a_1077_8251.n14 a_1077_8251.n43 18.7629
R2170 a_1077_8251.n43 a_1077_8251.n28 18.7629
R2171 a_1077_8251.n76 a_1077_8251.n75 27.1064
R2172 a_1077_8251.n45 a_1077_8251.n26 18.7629
R2173 a_1077_8251.n16 a_1077_8251.n47 18.7629
R2174 a_1077_8251.n47 a_1077_8251.n24 18.7629
R2175 a_1077_8251.n48 a_1077_8251.n3 18.7629
R2176 a_1077_8251.n49 a_1077_8251.n22 18.7629
R2177 a_1077_8251.n18 a_1077_8251.n51 18.7629
R2178 a_1077_8251.n51 a_1077_8251.n20 18.7629
R2179 a_1077_8251.n74 a_1077_8251.n11 33.5713
R2180 a_1077_8251.n7 a_1077_8251.t1 25.3133
R2181 a_1077_8251.n57 a_1077_8251.n53 13.2471
R2182 a_1077_8251.n58 a_1077_8251.n35 18.7629
R2183 a_1077_8251.n60 a_1077_8251.n33 18.7629
R2184 a_1077_8251.n61 a_1077_8251.n5 18.7629
R2185 a_1077_8251.n62 a_1077_8251.n31 18.7629
R2186 a_1077_8251.n64 a_1077_8251.n29 18.7629
R2187 a_1077_8251.n65 a_1077_8251.n55 13.2471
R2188 a_1077_8251.n66 a_1077_8251.n27 18.7629
R2189 a_1077_8251.n68 a_1077_8251.n25 18.7629
R2190 a_1077_8251.n69 a_1077_8251.n2 18.7629
R2191 a_1077_8251.n70 a_1077_8251.n23 18.7629
R2192 a_1077_8251.n72 a_1077_8251.n21 18.7629
R2193 a_1077_8251.n57 a_1077_8251.n35 18.7629
R2194 a_1077_8251.n58 a_1077_8251.n13 18.7629
R2195 a_1077_8251.n59 a_1077_8251.n33 18.7629
R2196 a_1077_8251.n60 a_1077_8251.n5 18.7629
R2197 a_1077_8251.n61 a_1077_8251.n31 18.7629
R2198 a_1077_8251.n62 a_1077_8251.n15 18.7629
R2199 a_1077_8251.n63 a_1077_8251.n29 18.7629
R2200 a_1077_8251.n64 a_1077_8251.n54 13.2471
R2201 a_1077_8251.n65 a_1077_8251.n27 18.7629
R2202 a_1077_8251.n66 a_1077_8251.n17 18.7629
R2203 a_1077_8251.n67 a_1077_8251.n25 18.7629
R2204 a_1077_8251.n68 a_1077_8251.n2 18.7629
R2205 a_1077_8251.n69 a_1077_8251.n23 18.7629
R2206 a_1077_8251.n70 a_1077_8251.n19 18.7629
R2207 a_1077_8251.n71 a_1077_8251.n21 18.7629
R2208 a_1077_8251.n72 a_1077_8251.n56 13.2471
R2209 a_1077_8251.n77 a_1077_8251.n37 13.2471
R2210 a_1077_8251.n75 a_1077_8251.n45 13.2471
R2211 a_1077_8251.n9 a_1077_8251.n36 53.1865
R2212 a_1077_8251.n76 a_1077_8251.n44 13.2471
R2213 a_1077_8251.n74 a_1077_8251.n52 13.2471
R2214 a_1077_8251.n7 a_1077_8251.n8 0.846729
R2215 a_1077_8251.n4 a_1077_8251.n53 9.3005
R2216 a_1077_8251.n4 a_1077_8251.n35 1.89332
R2217 a_1077_8251.n4 a_1077_8251.n13 1.89332
R2218 a_1077_8251.n4 a_1077_8251.n33 1.89332
R2219 a_1077_8251.n4 a_1077_8251.n5 1.89332
R2220 a_1077_8251.n4 a_1077_8251.n31 1.89332
R2221 a_1077_8251.n4 a_1077_8251.n15 1.89332
R2222 a_1077_8251.n4 a_1077_8251.n29 1.89332
R2223 a_1077_8251.n4 a_1077_8251.n54 9.3005
R2224 a_1077_8251.n1 a_1077_8251.n55 9.3005
R2225 a_1077_8251.n1 a_1077_8251.n27 1.89332
R2226 a_1077_8251.n1 a_1077_8251.n17 1.89332
R2227 a_1077_8251.n1 a_1077_8251.n25 1.89332
R2228 a_1077_8251.n1 a_1077_8251.n2 1.89332
R2229 a_1077_8251.n1 a_1077_8251.n23 1.89332
R2230 a_1077_8251.n1 a_1077_8251.n19 1.89332
R2231 a_1077_8251.n1 a_1077_8251.n21 1.89332
R2232 a_1077_8251.n1 a_1077_8251.n56 9.3005
R2233 a_1077_8251.n0 a_1077_8251.n10 0.77628
R2234 a_1077_8251.n10 a_1077_8251.n73 48.7551
R2235 a_1077_8251.n7 a_1077_8251.n9 0.846729
R2236 a_1077_8251.n9 a_1077_8251.n77 33.502
R2237 a_1077_8251.n77 a_1077_8251.n4 9.3005
R2238 a_1077_8251.n4 a_1077_8251.n34 1.89332
R2239 a_1077_8251.n38 a_1077_8251.n34 18.7629
R2240 a_1077_8251.n12 a_1077_8251.n38 18.7629
R2241 a_1077_8251.n12 a_1077_8251.n4 1.89332
R2242 a_1077_8251.n4 a_1077_8251.n32 1.89332
R2243 a_1077_8251.n40 a_1077_8251.n32 18.7629
R2244 a_1077_8251.n4 a_1077_8251.n6 1.89332
R2245 a_1077_8251.n41 a_1077_8251.n6 18.7629
R2246 a_1077_8251.n4 a_1077_8251.n30 1.89332
R2247 a_1077_8251.n42 a_1077_8251.n30 18.7629
R2248 a_1077_8251.n14 a_1077_8251.n42 18.7629
R2249 a_1077_8251.n14 a_1077_8251.n4 1.89332
R2250 a_1077_8251.n4 a_1077_8251.n28 1.89332
R2251 a_1077_8251.n44 a_1077_8251.n28 18.7629
R2252 a_1077_8251.n4 a_1077_8251.n76 9.3005
R2253 a_1077_8251.n75 a_1077_8251.n1 9.3005
R2254 a_1077_8251.n1 a_1077_8251.n26 1.89332
R2255 a_1077_8251.n46 a_1077_8251.n26 18.7629
R2256 a_1077_8251.n16 a_1077_8251.n46 18.7629
R2257 a_1077_8251.n16 a_1077_8251.n1 1.89332
R2258 a_1077_8251.n1 a_1077_8251.n24 1.89332
R2259 a_1077_8251.n48 a_1077_8251.n24 18.7629
R2260 a_1077_8251.n1 a_1077_8251.n3 1.89332
R2261 a_1077_8251.n49 a_1077_8251.n3 18.7629
R2262 a_1077_8251.n1 a_1077_8251.n22 1.89332
R2263 a_1077_8251.n50 a_1077_8251.n22 18.7629
R2264 a_1077_8251.n18 a_1077_8251.n50 18.7629
R2265 a_1077_8251.n18 a_1077_8251.n1 1.89332
R2266 a_1077_8251.n1 a_1077_8251.n20 1.89332
R2267 a_1077_8251.n52 a_1077_8251.n20 18.7629
R2268 a_1077_8251.n1 a_1077_8251.n74 9.3005
R2269 a_1077_8251.n11 a_1077_8251.n0 0.77628
R2270 a_1077_8251.n73 a_1077_8251.t2 1.433
R2271 a_1077_8251.t0 a_1077_8251.n36 1.433
R2272 a_1077_8251.n1 a_1077_8251.n0 0.336093
R2273 a_1077_8251.n7 a_1077_8251.n4 0.244568
R2274 a_1077_8251.n4 a_1077_8251.n1 0.244568
R2275 VDD.n1343 VDD.n1342 585
R2276 VDD.n256 VDD.n67 397.101
R2277 VDD.n259 VDD.n258 397.101
R2278 VDD.n217 VDD.n203 397.101
R2279 VDD.n249 VDD.n206 397.101
R2280 VDD.n169 VDD.n92 397.101
R2281 VDD.n171 VDD.n82 397.101
R2282 VDD.n130 VDD.n117 397.101
R2283 VDD.n162 VDD.n120 397.101
R2284 VDD.n803 VDD.n329 374.3
R2285 VDD.n813 VDD.n324 374.3
R2286 VDD.n792 VDD.n649 374.3
R2287 VDD.n795 VDD.n331 374.3
R2288 VDD.n635 VDD.n367 374.3
R2289 VDD.n645 VDD.n362 374.3
R2290 VDD.n519 VDD.n371 374.3
R2291 VDD.n522 VDD.n369 374.3
R2292 VDD.n1286 VDD.n945 355.3
R2293 VDD.n1330 VDD.n1329 355.3
R2294 VDD.n1298 VDD.n1297 355.3
R2295 VDD.n1291 VDD.n1290 355.3
R2296 VDD.n1122 VDD.n1121 355.3
R2297 VDD.n1012 VDD.n981 355.3
R2298 VDD.n1090 VDD.n1078 355.3
R2299 VDD.n1248 VDD.n975 355.3
R2300 VDD.n1339 VDD.t14 354.596
R2301 VDD.n1372 VDD.n1371 321.882
R2302 VDD.n1372 VDD.n40 321.882
R2303 VDD.n1376 VDD.n40 321.882
R2304 VDD.n1376 VDD.n34 321.882
R2305 VDD.n1394 VDD.n34 321.882
R2306 VDD.n1394 VDD.n31 321.882
R2307 VDD.n1398 VDD.n31 321.882
R2308 VDD.n1399 VDD.n1398 321.882
R2309 VDD.n1399 VDD.n3 321.882
R2310 VDD.n4 VDD.n3 321.882
R2311 VDD.n1404 VDD.n4 321.882
R2312 VDD.n1405 VDD.n1404 321.882
R2313 VDD.n1405 VDD.n9 321.882
R2314 VDD.n10 VDD.n9 321.882
R2315 VDD.n1409 VDD.n10 321.882
R2316 VDD.n1409 VDD.n13 321.882
R2317 VDD.n14 VDD.n13 321.882
R2318 VDD.n1413 VDD.n14 321.882
R2319 VDD.n1413 VDD.n18 321.882
R2320 VDD.n19 VDD.n18 321.882
R2321 VDD.n1417 VDD.n19 321.882
R2322 VDD.n1417 VDD.n23 321.882
R2323 VDD.n24 VDD.n23 321.882
R2324 VDD.n25 VDD.n24 321.882
R2325 VDD.n1422 VDD.n25 321.882
R2326 VDD.n1422 VDD.n29 321.882
R2327 VDD.n30 VDD.n29 321.882
R2328 VDD.n1370 VDD.n1369 318.757
R2329 VDD.n1426 VDD.n1425 318.757
R2330 VDD.n1343 VDD.n937 285.877
R2331 VDD.n1343 VDD.n936 285.877
R2332 VDD.n1343 VDD.n935 285.877
R2333 VDD.n1343 VDD.n934 285.877
R2334 VDD.n1343 VDD.n933 285.877
R2335 VDD.n1343 VDD.n932 285.877
R2336 VDD.n1343 VDD.n931 285.877
R2337 VDD.n1343 VDD.n930 285.877
R2338 VDD.n1343 VDD.n929 285.877
R2339 VDD.n1343 VDD.n928 285.877
R2340 VDD.n1344 VDD.n1343 285.877
R2341 VDD.n1343 VDD.n920 285.877
R2342 VDD.n1343 VDD.n919 285.877
R2343 VDD.n1460 VDD.t33 257.618
R2344 VDD.n1 VDD.t1 257.618
R2345 VDD.n1429 VDD.t23 249.873
R2346 VDD.n1366 VDD.t8 249.873
R2347 VDD.n1466 VDD.t37 249.873
R2348 VDD.n1453 VDD.t20 249.873
R2349 VDD.n1286 VDD.n1285 185
R2350 VDD.n1284 VDD.n1257 185
R2351 VDD.n1283 VDD.n1256 185
R2352 VDD.n1288 VDD.n1256 185
R2353 VDD.n1282 VDD.n1281 185
R2354 VDD.n1280 VDD.n1279 185
R2355 VDD.n1278 VDD.n1277 185
R2356 VDD.n1276 VDD.n1275 185
R2357 VDD.n1274 VDD.n1273 185
R2358 VDD.n1272 VDD.n1271 185
R2359 VDD.n1270 VDD.n1269 185
R2360 VDD.n1268 VDD.n1267 185
R2361 VDD.n1266 VDD.n1265 185
R2362 VDD.n1264 VDD.n1263 185
R2363 VDD.n1262 VDD.n1261 185
R2364 VDD.n1260 VDD.n1259 185
R2365 VDD.n1258 VDD.n964 185
R2366 VDD.n1290 VDD.n963 185
R2367 VDD.n1299 VDD.n1298 185
R2368 VDD.n1301 VDD.n1300 185
R2369 VDD.n1303 VDD.n1302 185
R2370 VDD.n1305 VDD.n1304 185
R2371 VDD.n1307 VDD.n1306 185
R2372 VDD.n1309 VDD.n1308 185
R2373 VDD.n1311 VDD.n1310 185
R2374 VDD.n1313 VDD.n1312 185
R2375 VDD.n1315 VDD.n1314 185
R2376 VDD.n1317 VDD.n1316 185
R2377 VDD.n1319 VDD.n1318 185
R2378 VDD.n1321 VDD.n1320 185
R2379 VDD.n1323 VDD.n1322 185
R2380 VDD.n1324 VDD.n961 185
R2381 VDD.n1326 VDD.n1325 185
R2382 VDD.n962 VDD.n952 185
R2383 VDD.n1329 VDD.n953 185
R2384 VDD.n1329 VDD.n1328 185
R2385 VDD.n1297 VDD.n1296 185
R2386 VDD.n1297 VDD.n951 185
R2387 VDD.n1295 VDD.n950 185
R2388 VDD.n1333 VDD.n950 185
R2389 VDD.n1294 VDD.n949 185
R2390 VDD.n1334 VDD.n949 185
R2391 VDD.n1293 VDD.n948 185
R2392 VDD.n1335 VDD.n948 185
R2393 VDD.n1292 VDD.n1291 185
R2394 VDD.n1291 VDD.n947 185
R2395 VDD.n945 VDD.n943 185
R2396 VDD.n947 VDD.n945 185
R2397 VDD.n1337 VDD.n1336 185
R2398 VDD.n1336 VDD.n1335 185
R2399 VDD.n946 VDD.n944 185
R2400 VDD.n1334 VDD.n946 185
R2401 VDD.n1332 VDD.n1331 185
R2402 VDD.n1333 VDD.n1332 185
R2403 VDD.n1330 VDD.n941 185
R2404 VDD.n1330 VDD.n951 185
R2405 VDD.n1248 VDD.n1247 185
R2406 VDD.n1249 VDD.n1248 185
R2407 VDD.n976 VDD.n974 185
R2408 VDD.n983 VDD.n982 185
R2409 VDD.n985 VDD.n984 185
R2410 VDD.n987 VDD.n986 185
R2411 VDD.n989 VDD.n988 185
R2412 VDD.n991 VDD.n990 185
R2413 VDD.n993 VDD.n992 185
R2414 VDD.n995 VDD.n994 185
R2415 VDD.n997 VDD.n996 185
R2416 VDD.n999 VDD.n998 185
R2417 VDD.n1001 VDD.n1000 185
R2418 VDD.n1003 VDD.n1002 185
R2419 VDD.n1005 VDD.n1004 185
R2420 VDD.n1007 VDD.n1006 185
R2421 VDD.n1009 VDD.n1008 185
R2422 VDD.n1010 VDD.n981 185
R2423 VDD.n1246 VDD.n975 185
R2424 VDD.n975 VDD.n965 185
R2425 VDD.n1245 VDD.n1244 185
R2426 VDD.n1244 VDD.n1243 185
R2427 VDD.n978 VDD.n977 185
R2428 VDD.n979 VDD.n978 185
R2429 VDD.n1226 VDD.n1225 185
R2430 VDD.n1227 VDD.n1226 185
R2431 VDD.n1224 VDD.n1022 185
R2432 VDD.n1228 VDD.n1022 185
R2433 VDD.n1223 VDD.n1021 185
R2434 VDD.n1229 VDD.n1021 185
R2435 VDD.n1222 VDD.n1221 185
R2436 VDD.n1221 VDD.n1020 185
R2437 VDD.n1220 VDD.n1023 185
R2438 VDD.n1220 VDD.n1219 185
R2439 VDD.n1201 VDD.n1024 185
R2440 VDD.n1025 VDD.n1024 185
R2441 VDD.n1203 VDD.n1202 185
R2442 VDD.n1204 VDD.n1203 185
R2443 VDD.n1200 VDD.n1033 185
R2444 VDD.n1033 VDD.n1032 185
R2445 VDD.n1199 VDD.n1198 185
R2446 VDD.n1198 VDD.n1197 185
R2447 VDD.n1035 VDD.n1034 185
R2448 VDD.n1036 VDD.n1035 185
R2449 VDD.n1181 VDD.n1180 185
R2450 VDD.n1182 VDD.n1181 185
R2451 VDD.n1179 VDD.n1044 185
R2452 VDD.n1044 VDD.n1043 185
R2453 VDD.n1178 VDD.n1177 185
R2454 VDD.n1177 VDD.n1176 185
R2455 VDD.n1046 VDD.n1045 185
R2456 VDD.n1047 VDD.n1046 185
R2457 VDD.n1160 VDD.n1159 185
R2458 VDD.n1161 VDD.n1160 185
R2459 VDD.n1158 VDD.n1055 185
R2460 VDD.n1055 VDD.n1054 185
R2461 VDD.n1157 VDD.n1156 185
R2462 VDD.n1156 VDD.n1155 185
R2463 VDD.n1057 VDD.n1056 185
R2464 VDD.n1058 VDD.n1057 185
R2465 VDD.n1139 VDD.n1138 185
R2466 VDD.n1140 VDD.n1139 185
R2467 VDD.n1137 VDD.n1069 185
R2468 VDD.n1069 VDD.n1068 185
R2469 VDD.n1136 VDD.n1135 185
R2470 VDD.n1135 VDD.n1134 185
R2471 VDD.n1071 VDD.n1070 185
R2472 VDD.n1132 VDD.n1071 185
R2473 VDD.n1130 VDD.n1129 185
R2474 VDD.n1131 VDD.n1130 185
R2475 VDD.n1128 VDD.n1074 185
R2476 VDD.n1074 VDD.n1073 185
R2477 VDD.n1127 VDD.n1126 185
R2478 VDD.n1126 VDD.n1125 185
R2479 VDD.n1076 VDD.n1075 185
R2480 VDD.n1124 VDD.n1076 185
R2481 VDD.n1088 VDD.n1078 185
R2482 VDD.n1123 VDD.n1078 185
R2483 VDD.n1121 VDD.n1120 185
R2484 VDD.n1119 VDD.n1118 185
R2485 VDD.n1117 VDD.n1080 185
R2486 VDD.n1117 VDD.n1077 185
R2487 VDD.n1116 VDD.n1115 185
R2488 VDD.n1114 VDD.n1113 185
R2489 VDD.n1112 VDD.n1082 185
R2490 VDD.n1110 VDD.n1109 185
R2491 VDD.n1108 VDD.n1083 185
R2492 VDD.n1107 VDD.n1106 185
R2493 VDD.n1104 VDD.n1084 185
R2494 VDD.n1102 VDD.n1101 185
R2495 VDD.n1100 VDD.n1085 185
R2496 VDD.n1099 VDD.n1098 185
R2497 VDD.n1096 VDD.n1086 185
R2498 VDD.n1094 VDD.n1093 185
R2499 VDD.n1092 VDD.n1087 185
R2500 VDD.n1091 VDD.n1090 185
R2501 VDD.n1012 VDD.n1011 185
R2502 VDD.n1012 VDD.n965 185
R2503 VDD.n1242 VDD.n1241 185
R2504 VDD.n1243 VDD.n1242 185
R2505 VDD.n1240 VDD.n980 185
R2506 VDD.n980 VDD.n979 185
R2507 VDD.n1239 VDD.n1014 185
R2508 VDD.n1227 VDD.n1014 185
R2509 VDD.n1019 VDD.n1013 185
R2510 VDD.n1228 VDD.n1019 185
R2511 VDD.n1231 VDD.n1230 185
R2512 VDD.n1230 VDD.n1229 185
R2513 VDD.n1018 VDD.n1017 185
R2514 VDD.n1020 VDD.n1018 185
R2515 VDD.n1218 VDD.n1217 185
R2516 VDD.n1219 VDD.n1218 185
R2517 VDD.n1027 VDD.n1026 185
R2518 VDD.n1026 VDD.n1025 185
R2519 VDD.n1206 VDD.n1205 185
R2520 VDD.n1205 VDD.n1204 185
R2521 VDD.n1031 VDD.n1030 185
R2522 VDD.n1032 VDD.n1031 185
R2523 VDD.n1196 VDD.n1195 185
R2524 VDD.n1197 VDD.n1196 185
R2525 VDD.n1038 VDD.n1037 185
R2526 VDD.n1037 VDD.n1036 185
R2527 VDD.n1184 VDD.n1183 185
R2528 VDD.n1183 VDD.n1182 185
R2529 VDD.n1042 VDD.n1041 185
R2530 VDD.n1043 VDD.n1042 185
R2531 VDD.n1175 VDD.n1174 185
R2532 VDD.n1176 VDD.n1175 185
R2533 VDD.n1049 VDD.n1048 185
R2534 VDD.n1048 VDD.n1047 185
R2535 VDD.n1163 VDD.n1162 185
R2536 VDD.n1162 VDD.n1161 185
R2537 VDD.n1053 VDD.n1052 185
R2538 VDD.n1054 VDD.n1053 185
R2539 VDD.n1154 VDD.n1153 185
R2540 VDD.n1155 VDD.n1154 185
R2541 VDD.n1060 VDD.n1059 185
R2542 VDD.n1059 VDD.n1058 185
R2543 VDD.n1142 VDD.n1141 185
R2544 VDD.n1141 VDD.n1140 185
R2545 VDD.n1067 VDD.n1066 185
R2546 VDD.n1068 VDD.n1067 185
R2547 VDD.n1133 VDD.n924 185
R2548 VDD.n1134 VDD.n1133 185
R2549 VDD.n1348 VDD.n923 185
R2550 VDD.n1132 VDD.n923 185
R2551 VDD.n1349 VDD.n922 185
R2552 VDD.n1131 VDD.n922 185
R2553 VDD.n1072 VDD.n917 185
R2554 VDD.n1073 VDD.n1072 185
R2555 VDD.n1356 VDD.n916 185
R2556 VDD.n1125 VDD.n916 185
R2557 VDD.n1357 VDD.n915 185
R2558 VDD.n1124 VDD.n915 185
R2559 VDD.n1122 VDD.n913 185
R2560 VDD.n1123 VDD.n1122 185
R2561 VDD.n805 VDD.n329 185
R2562 VDD.n329 VDD.n327 185
R2563 VDD.n807 VDD.n806 185
R2564 VDD.n808 VDD.n807 185
R2565 VDD.n797 VDD.n328 185
R2566 VDD.n793 VDD.n328 185
R2567 VDD.n796 VDD.n795 185
R2568 VDD.n795 VDD.n794 185
R2569 VDD.n331 VDD.n330 185
R2570 VDD.n680 VDD.n678 185
R2571 VDD.n681 VDD.n677 185
R2572 VDD.n681 VDD.n648 185
R2573 VDD.n684 VDD.n683 185
R2574 VDD.n685 VDD.n676 185
R2575 VDD.n687 VDD.n686 185
R2576 VDD.n689 VDD.n675 185
R2577 VDD.n692 VDD.n691 185
R2578 VDD.n693 VDD.n674 185
R2579 VDD.n695 VDD.n694 185
R2580 VDD.n697 VDD.n673 185
R2581 VDD.n700 VDD.n699 185
R2582 VDD.n701 VDD.n672 185
R2583 VDD.n703 VDD.n702 185
R2584 VDD.n705 VDD.n671 185
R2585 VDD.n708 VDD.n707 185
R2586 VDD.n709 VDD.n670 185
R2587 VDD.n711 VDD.n710 185
R2588 VDD.n713 VDD.n669 185
R2589 VDD.n716 VDD.n715 185
R2590 VDD.n717 VDD.n668 185
R2591 VDD.n719 VDD.n718 185
R2592 VDD.n721 VDD.n667 185
R2593 VDD.n724 VDD.n723 185
R2594 VDD.n725 VDD.n666 185
R2595 VDD.n727 VDD.n726 185
R2596 VDD.n729 VDD.n665 185
R2597 VDD.n732 VDD.n731 185
R2598 VDD.n733 VDD.n664 185
R2599 VDD.n735 VDD.n734 185
R2600 VDD.n737 VDD.n663 185
R2601 VDD.n740 VDD.n739 185
R2602 VDD.n741 VDD.n662 185
R2603 VDD.n743 VDD.n742 185
R2604 VDD.n745 VDD.n661 185
R2605 VDD.n748 VDD.n747 185
R2606 VDD.n749 VDD.n660 185
R2607 VDD.n751 VDD.n750 185
R2608 VDD.n753 VDD.n659 185
R2609 VDD.n756 VDD.n755 185
R2610 VDD.n757 VDD.n658 185
R2611 VDD.n759 VDD.n758 185
R2612 VDD.n761 VDD.n657 185
R2613 VDD.n764 VDD.n763 185
R2614 VDD.n765 VDD.n656 185
R2615 VDD.n767 VDD.n766 185
R2616 VDD.n769 VDD.n655 185
R2617 VDD.n772 VDD.n771 185
R2618 VDD.n773 VDD.n654 185
R2619 VDD.n775 VDD.n774 185
R2620 VDD.n777 VDD.n653 185
R2621 VDD.n780 VDD.n779 185
R2622 VDD.n781 VDD.n652 185
R2623 VDD.n783 VDD.n782 185
R2624 VDD.n785 VDD.n651 185
R2625 VDD.n786 VDD.n650 185
R2626 VDD.n789 VDD.n788 185
R2627 VDD.n790 VDD.n649 185
R2628 VDD.n649 VDD.n648 185
R2629 VDD.n813 VDD.n812 185
R2630 VDD.n815 VDD.n322 185
R2631 VDD.n817 VDD.n816 185
R2632 VDD.n818 VDD.n321 185
R2633 VDD.n820 VDD.n819 185
R2634 VDD.n822 VDD.n319 185
R2635 VDD.n824 VDD.n823 185
R2636 VDD.n825 VDD.n318 185
R2637 VDD.n827 VDD.n826 185
R2638 VDD.n829 VDD.n316 185
R2639 VDD.n831 VDD.n830 185
R2640 VDD.n832 VDD.n315 185
R2641 VDD.n834 VDD.n833 185
R2642 VDD.n836 VDD.n313 185
R2643 VDD.n838 VDD.n837 185
R2644 VDD.n839 VDD.n312 185
R2645 VDD.n841 VDD.n840 185
R2646 VDD.n843 VDD.n310 185
R2647 VDD.n845 VDD.n844 185
R2648 VDD.n846 VDD.n309 185
R2649 VDD.n848 VDD.n847 185
R2650 VDD.n850 VDD.n307 185
R2651 VDD.n852 VDD.n851 185
R2652 VDD.n853 VDD.n306 185
R2653 VDD.n855 VDD.n854 185
R2654 VDD.n857 VDD.n304 185
R2655 VDD.n859 VDD.n858 185
R2656 VDD.n860 VDD.n303 185
R2657 VDD.n862 VDD.n861 185
R2658 VDD.n864 VDD.n301 185
R2659 VDD.n866 VDD.n865 185
R2660 VDD.n867 VDD.n300 185
R2661 VDD.n869 VDD.n868 185
R2662 VDD.n871 VDD.n298 185
R2663 VDD.n873 VDD.n872 185
R2664 VDD.n874 VDD.n297 185
R2665 VDD.n876 VDD.n875 185
R2666 VDD.n878 VDD.n295 185
R2667 VDD.n880 VDD.n879 185
R2668 VDD.n881 VDD.n294 185
R2669 VDD.n883 VDD.n882 185
R2670 VDD.n885 VDD.n292 185
R2671 VDD.n887 VDD.n886 185
R2672 VDD.n888 VDD.n291 185
R2673 VDD.n890 VDD.n889 185
R2674 VDD.n892 VDD.n289 185
R2675 VDD.n894 VDD.n893 185
R2676 VDD.n895 VDD.n288 185
R2677 VDD.n897 VDD.n896 185
R2678 VDD.n899 VDD.n286 185
R2679 VDD.n901 VDD.n900 185
R2680 VDD.n903 VDD.n284 185
R2681 VDD.n905 VDD.n904 185
R2682 VDD.n907 VDD.n281 185
R2683 VDD.n909 VDD.n908 185
R2684 VDD.n799 VDD.n280 185
R2685 VDD.n801 VDD.n800 185
R2686 VDD.n804 VDD.n803 185
R2687 VDD.n811 VDD.n324 185
R2688 VDD.n327 VDD.n324 185
R2689 VDD.n810 VDD.n809 185
R2690 VDD.n809 VDD.n808 185
R2691 VDD.n326 VDD.n325 185
R2692 VDD.n793 VDD.n326 185
R2693 VDD.n792 VDD.n791 185
R2694 VDD.n794 VDD.n792 185
R2695 VDD.n637 VDD.n367 185
R2696 VDD.n367 VDD.n332 185
R2697 VDD.n639 VDD.n638 185
R2698 VDD.n640 VDD.n639 185
R2699 VDD.n524 VDD.n366 185
R2700 VDD.n520 VDD.n366 185
R2701 VDD.n523 VDD.n522 185
R2702 VDD.n522 VDD.n521 185
R2703 VDD.n645 VDD.n644 185
R2704 VDD.n363 VDD.n361 185
R2705 VDD.n526 VDD.n525 185
R2706 VDD.n528 VDD.n527 185
R2707 VDD.n530 VDD.n529 185
R2708 VDD.n532 VDD.n531 185
R2709 VDD.n534 VDD.n533 185
R2710 VDD.n536 VDD.n535 185
R2711 VDD.n538 VDD.n537 185
R2712 VDD.n540 VDD.n539 185
R2713 VDD.n542 VDD.n541 185
R2714 VDD.n544 VDD.n543 185
R2715 VDD.n546 VDD.n545 185
R2716 VDD.n548 VDD.n547 185
R2717 VDD.n550 VDD.n549 185
R2718 VDD.n552 VDD.n551 185
R2719 VDD.n554 VDD.n553 185
R2720 VDD.n556 VDD.n555 185
R2721 VDD.n558 VDD.n557 185
R2722 VDD.n560 VDD.n559 185
R2723 VDD.n562 VDD.n561 185
R2724 VDD.n564 VDD.n563 185
R2725 VDD.n566 VDD.n565 185
R2726 VDD.n568 VDD.n567 185
R2727 VDD.n570 VDD.n569 185
R2728 VDD.n572 VDD.n571 185
R2729 VDD.n574 VDD.n573 185
R2730 VDD.n576 VDD.n575 185
R2731 VDD.n578 VDD.n577 185
R2732 VDD.n580 VDD.n579 185
R2733 VDD.n582 VDD.n581 185
R2734 VDD.n584 VDD.n583 185
R2735 VDD.n586 VDD.n585 185
R2736 VDD.n588 VDD.n587 185
R2737 VDD.n590 VDD.n589 185
R2738 VDD.n592 VDD.n591 185
R2739 VDD.n594 VDD.n593 185
R2740 VDD.n596 VDD.n595 185
R2741 VDD.n598 VDD.n597 185
R2742 VDD.n600 VDD.n599 185
R2743 VDD.n602 VDD.n601 185
R2744 VDD.n604 VDD.n603 185
R2745 VDD.n606 VDD.n605 185
R2746 VDD.n608 VDD.n607 185
R2747 VDD.n610 VDD.n609 185
R2748 VDD.n612 VDD.n611 185
R2749 VDD.n614 VDD.n613 185
R2750 VDD.n616 VDD.n615 185
R2751 VDD.n618 VDD.n617 185
R2752 VDD.n620 VDD.n619 185
R2753 VDD.n622 VDD.n621 185
R2754 VDD.n624 VDD.n623 185
R2755 VDD.n626 VDD.n625 185
R2756 VDD.n628 VDD.n627 185
R2757 VDD.n630 VDD.n629 185
R2758 VDD.n632 VDD.n631 185
R2759 VDD.n634 VDD.n633 185
R2760 VDD.n636 VDD.n635 185
R2761 VDD.n643 VDD.n362 185
R2762 VDD.n362 VDD.n332 185
R2763 VDD.n642 VDD.n641 185
R2764 VDD.n641 VDD.n640 185
R2765 VDD.n365 VDD.n364 185
R2766 VDD.n520 VDD.n365 185
R2767 VDD.n519 VDD.n518 185
R2768 VDD.n521 VDD.n519 185
R2769 VDD.n369 VDD.n368 185
R2770 VDD.n405 VDD.n403 185
R2771 VDD.n406 VDD.n400 185
R2772 VDD.n406 VDD.n370 185
R2773 VDD.n409 VDD.n408 185
R2774 VDD.n410 VDD.n399 185
R2775 VDD.n414 VDD.n413 185
R2776 VDD.n416 VDD.n398 185
R2777 VDD.n419 VDD.n418 185
R2778 VDD.n420 VDD.n396 185
R2779 VDD.n422 VDD.n421 185
R2780 VDD.n424 VDD.n395 185
R2781 VDD.n427 VDD.n426 185
R2782 VDD.n428 VDD.n394 185
R2783 VDD.n430 VDD.n429 185
R2784 VDD.n432 VDD.n393 185
R2785 VDD.n435 VDD.n434 185
R2786 VDD.n436 VDD.n392 185
R2787 VDD.n438 VDD.n437 185
R2788 VDD.n440 VDD.n391 185
R2789 VDD.n443 VDD.n442 185
R2790 VDD.n444 VDD.n390 185
R2791 VDD.n446 VDD.n445 185
R2792 VDD.n448 VDD.n389 185
R2793 VDD.n451 VDD.n450 185
R2794 VDD.n452 VDD.n388 185
R2795 VDD.n454 VDD.n453 185
R2796 VDD.n456 VDD.n387 185
R2797 VDD.n459 VDD.n458 185
R2798 VDD.n460 VDD.n386 185
R2799 VDD.n462 VDD.n461 185
R2800 VDD.n464 VDD.n385 185
R2801 VDD.n467 VDD.n466 185
R2802 VDD.n468 VDD.n384 185
R2803 VDD.n470 VDD.n469 185
R2804 VDD.n472 VDD.n383 185
R2805 VDD.n475 VDD.n474 185
R2806 VDD.n476 VDD.n382 185
R2807 VDD.n478 VDD.n477 185
R2808 VDD.n480 VDD.n381 185
R2809 VDD.n483 VDD.n482 185
R2810 VDD.n484 VDD.n380 185
R2811 VDD.n486 VDD.n485 185
R2812 VDD.n488 VDD.n379 185
R2813 VDD.n491 VDD.n490 185
R2814 VDD.n492 VDD.n378 185
R2815 VDD.n494 VDD.n493 185
R2816 VDD.n496 VDD.n377 185
R2817 VDD.n499 VDD.n498 185
R2818 VDD.n500 VDD.n376 185
R2819 VDD.n502 VDD.n501 185
R2820 VDD.n504 VDD.n375 185
R2821 VDD.n507 VDD.n506 185
R2822 VDD.n508 VDD.n374 185
R2823 VDD.n510 VDD.n509 185
R2824 VDD.n512 VDD.n373 185
R2825 VDD.n513 VDD.n372 185
R2826 VDD.n516 VDD.n515 185
R2827 VDD.n517 VDD.n371 185
R2828 VDD.n371 VDD.n370 185
R2829 VDD.n249 VDD.n248 185
R2830 VDD.n250 VDD.n249 185
R2831 VDD.n208 VDD.n204 185
R2832 VDD.n251 VDD.n204 185
R2833 VDD.n207 VDD.n64 185
R2834 VDD.n66 VDD.n64 185
R2835 VDD.n258 VDD.n65 185
R2836 VDD.n258 VDD.n257 185
R2837 VDD.n247 VDD.n206 185
R2838 VDD.n246 VDD.n245 185
R2839 VDD.n243 VDD.n209 185
R2840 VDD.n241 VDD.n240 185
R2841 VDD.n239 VDD.n210 185
R2842 VDD.n238 VDD.n237 185
R2843 VDD.n235 VDD.n211 185
R2844 VDD.n233 VDD.n232 185
R2845 VDD.n231 VDD.n212 185
R2846 VDD.n230 VDD.n229 185
R2847 VDD.n227 VDD.n213 185
R2848 VDD.n225 VDD.n224 185
R2849 VDD.n223 VDD.n214 185
R2850 VDD.n222 VDD.n221 185
R2851 VDD.n219 VDD.n215 185
R2852 VDD.n217 VDD.n216 185
R2853 VDD.n256 VDD.n255 185
R2854 VDD.n257 VDD.n256 185
R2855 VDD.n254 VDD.n68 185
R2856 VDD.n68 VDD.n66 185
R2857 VDD.n253 VDD.n252 185
R2858 VDD.n252 VDD.n251 185
R2859 VDD.n203 VDD.n202 185
R2860 VDD.n250 VDD.n203 185
R2861 VDD.n259 VDD.n56 185
R2862 VDD.n262 VDD.n261 185
R2863 VDD.n57 VDD.n55 185
R2864 VDD.n266 VDD.n54 185
R2865 VDD.n267 VDD.n53 185
R2866 VDD.n268 VDD.n52 185
R2867 VDD.n59 VDD.n49 185
R2868 VDD.n272 VDD.n48 185
R2869 VDD.n273 VDD.n47 185
R2870 VDD.n274 VDD.n46 185
R2871 VDD.n191 VDD.n45 185
R2872 VDD.n195 VDD.n193 185
R2873 VDD.n196 VDD.n190 185
R2874 VDD.n197 VDD.n188 185
R2875 VDD.n187 VDD.n69 185
R2876 VDD.n201 VDD.n67 185
R2877 VDD.n162 VDD.n161 185
R2878 VDD.n163 VDD.n162 185
R2879 VDD.n121 VDD.n118 185
R2880 VDD.n164 VDD.n118 185
R2881 VDD.n84 VDD.n83 185
R2882 VDD.n91 VDD.n84 185
R2883 VDD.n172 VDD.n171 185
R2884 VDD.n171 VDD.n170 185
R2885 VDD.n160 VDD.n120 185
R2886 VDD.n159 VDD.n158 185
R2887 VDD.n156 VDD.n122 185
R2888 VDD.n154 VDD.n153 185
R2889 VDD.n152 VDD.n123 185
R2890 VDD.n151 VDD.n150 185
R2891 VDD.n148 VDD.n124 185
R2892 VDD.n146 VDD.n145 185
R2893 VDD.n144 VDD.n125 185
R2894 VDD.n143 VDD.n142 185
R2895 VDD.n140 VDD.n126 185
R2896 VDD.n138 VDD.n137 185
R2897 VDD.n136 VDD.n127 185
R2898 VDD.n135 VDD.n134 185
R2899 VDD.n132 VDD.n128 185
R2900 VDD.n130 VDD.n129 185
R2901 VDD.n169 VDD.n168 185
R2902 VDD.n170 VDD.n169 185
R2903 VDD.n167 VDD.n93 185
R2904 VDD.n93 VDD.n91 185
R2905 VDD.n166 VDD.n165 185
R2906 VDD.n165 VDD.n164 185
R2907 VDD.n117 VDD.n116 185
R2908 VDD.n163 VDD.n117 185
R2909 VDD.n173 VDD.n82 185
R2910 VDD.n175 VDD.n81 185
R2911 VDD.n176 VDD.n80 185
R2912 VDD.n177 VDD.n79 185
R2913 VDD.n86 VDD.n77 185
R2914 VDD.n181 VDD.n76 185
R2915 VDD.n182 VDD.n75 185
R2916 VDD.n183 VDD.n74 185
R2917 VDD.n104 VDD.n73 185
R2918 VDD.n107 VDD.n106 185
R2919 VDD.n108 VDD.n103 185
R2920 VDD.n110 VDD.n101 185
R2921 VDD.n111 VDD.n100 185
R2922 VDD.n112 VDD.n98 185
R2923 VDD.n97 VDD.n94 185
R2924 VDD.n115 VDD.n92 185
R2925 VDD.n1432 VDD.n30 185
R2926 VDD.n1433 VDD.n29 185
R2927 VDD.n1424 VDD.n29 185
R2928 VDD.n1422 VDD.n26 185
R2929 VDD.n1423 VDD.n1422 185
R2930 VDD.n1440 VDD.n25 185
R2931 VDD.n1421 VDD.n25 185
R2932 VDD.n1441 VDD.n24 185
R2933 VDD.n1420 VDD.n24 185
R2934 VDD.n1442 VDD.n23 185
R2935 VDD.n1419 VDD.n23 185
R2936 VDD.n1417 VDD.n20 185
R2937 VDD.n1418 VDD.n1417 185
R2938 VDD.n1449 VDD.n19 185
R2939 VDD.n1416 VDD.n19 185
R2940 VDD.n1450 VDD.n18 185
R2941 VDD.n1415 VDD.n18 185
R2942 VDD.n1413 VDD.n15 185
R2943 VDD.n1414 VDD.n1413 185
R2944 VDD.n1456 VDD.n14 185
R2945 VDD.n1412 VDD.n14 185
R2946 VDD.n1457 VDD.n13 185
R2947 VDD.n1411 VDD.n13 185
R2948 VDD.n1409 VDD.n11 185
R2949 VDD.n1410 VDD.n1409 185
R2950 VDD.n1462 VDD.n10 185
R2951 VDD.n1408 VDD.n10 185
R2952 VDD.n1463 VDD.n9 185
R2953 VDD.n1407 VDD.n9 185
R2954 VDD.n1405 VDD.n8 185
R2955 VDD.n1406 VDD.n1405 185
R2956 VDD.n1404 VDD.n5 185
R2957 VDD.n1404 VDD.n1403 185
R2958 VDD.n1470 VDD.n4 185
R2959 VDD.n1402 VDD.n4 185
R2960 VDD.n1471 VDD.n3 185
R2961 VDD.n1401 VDD.n3 185
R2962 VDD.n1399 VDD.n2 185
R2963 VDD.n1400 VDD.n1399 185
R2964 VDD.n1398 VDD.n32 185
R2965 VDD.n1398 VDD.n1397 185
R2966 VDD.n36 VDD.n31 185
R2967 VDD.n1396 VDD.n31 185
R2968 VDD.n1394 VDD.n1393 185
R2969 VDD.n1395 VDD.n1394 185
R2970 VDD.n35 VDD.n34 185
R2971 VDD.n34 VDD.n33 185
R2972 VDD.n1377 VDD.n1376 185
R2973 VDD.n1376 VDD.n1375 185
R2974 VDD.n1378 VDD.n40 185
R2975 VDD.n1374 VDD.n40 185
R2976 VDD.n1372 VDD.n39 185
R2977 VDD.n1373 VDD.n1372 185
R2978 VDD.n1371 VDD.n41 185
R2979 VDD.n1370 VDD.t7 177.357
R2980 VDD.n1425 VDD.t22 177.357
R2981 VDD.n1374 VDD.n1373 175.386
R2982 VDD.n1395 VDD.n33 175.386
R2983 VDD.n1397 VDD.n1396 175.386
R2984 VDD.n1401 VDD.n1400 175.386
R2985 VDD.n1403 VDD.n1402 175.386
R2986 VDD.n1407 VDD.n1406 175.386
R2987 VDD.n1408 VDD.n1407 175.386
R2988 VDD.n1411 VDD.n1410 175.386
R2989 VDD.n1414 VDD.n1412 175.386
R2990 VDD.n1415 VDD.n1414 175.386
R2991 VDD.n1418 VDD.n1416 175.386
R2992 VDD.n1420 VDD.n1419 175.386
R2993 VDD.n1424 VDD.n1423 175.386
R2994 VDD.t0 VDD.n1401 169.905
R2995 VDD.t32 VDD.n1408 169.905
R2996 VDD.n1400 VDD.t30 162.596
R2997 VDD.t34 VDD.n1415 162.596
R2998 VDD.n1437 VDD.n1436 151.093
R2999 VDD.n1382 VDD.n1381 151.093
R3000 VDD.n1390 VDD.n1387 150.921
R3001 VDD.n1446 VDD.n1445 150.921
R3002 VDD.n1288 VDD.n1249 145.698
R3003 VDD.n1375 VDD.t9 144.327
R3004 VDD.n1421 VDD.t28 144.327
R3005 VDD.n1375 VDD.t11 140.673
R3006 VDD.t24 VDD.n1421 140.673
R3007 VDD.n1336 VDD.n945 136.8
R3008 VDD.n1336 VDD.n946 136.8
R3009 VDD.n1332 VDD.n946 136.8
R3010 VDD.n1332 VDD.n1330 136.8
R3011 VDD.n1329 VDD.n952 136.8
R3012 VDD.n1326 VDD.n961 136.8
R3013 VDD.n1322 VDD.n1321 136.8
R3014 VDD.n1318 VDD.n1317 136.8
R3015 VDD.n1314 VDD.n1313 136.8
R3016 VDD.n1310 VDD.n1309 136.8
R3017 VDD.n1306 VDD.n1305 136.8
R3018 VDD.n1302 VDD.n1301 136.8
R3019 VDD.n1291 VDD.n948 136.8
R3020 VDD.n949 VDD.n948 136.8
R3021 VDD.n950 VDD.n949 136.8
R3022 VDD.n1297 VDD.n950 136.8
R3023 VDD.n1257 VDD.n1256 136.8
R3024 VDD.n1281 VDD.n1256 136.8
R3025 VDD.n1279 VDD.n1278 136.8
R3026 VDD.n1275 VDD.n1274 136.8
R3027 VDD.n1271 VDD.n1270 136.8
R3028 VDD.n1267 VDD.n1266 136.8
R3029 VDD.n1263 VDD.n1262 136.8
R3030 VDD.n1259 VDD.n964 136.8
R3031 VDD.n1122 VDD.n915 136.8
R3032 VDD.n916 VDD.n915 136.8
R3033 VDD.n1072 VDD.n916 136.8
R3034 VDD.n1072 VDD.n922 136.8
R3035 VDD.n923 VDD.n922 136.8
R3036 VDD.n1133 VDD.n923 136.8
R3037 VDD.n1133 VDD.n1067 136.8
R3038 VDD.n1141 VDD.n1067 136.8
R3039 VDD.n1141 VDD.n1059 136.8
R3040 VDD.n1154 VDD.n1059 136.8
R3041 VDD.n1154 VDD.n1053 136.8
R3042 VDD.n1162 VDD.n1053 136.8
R3043 VDD.n1162 VDD.n1048 136.8
R3044 VDD.n1175 VDD.n1048 136.8
R3045 VDD.n1175 VDD.n1042 136.8
R3046 VDD.n1183 VDD.n1042 136.8
R3047 VDD.n1183 VDD.n1037 136.8
R3048 VDD.n1196 VDD.n1037 136.8
R3049 VDD.n1196 VDD.n1031 136.8
R3050 VDD.n1205 VDD.n1031 136.8
R3051 VDD.n1205 VDD.n1026 136.8
R3052 VDD.n1218 VDD.n1026 136.8
R3053 VDD.n1218 VDD.n1018 136.8
R3054 VDD.n1230 VDD.n1018 136.8
R3055 VDD.n1230 VDD.n1019 136.8
R3056 VDD.n1019 VDD.n1014 136.8
R3057 VDD.n1014 VDD.n980 136.8
R3058 VDD.n1242 VDD.n980 136.8
R3059 VDD.n1242 VDD.n1012 136.8
R3060 VDD.n1118 VDD.n1117 136.8
R3061 VDD.n1117 VDD.n1116 136.8
R3062 VDD.n1113 VDD.n1112 136.8
R3063 VDD.n1110 VDD.n1083 136.8
R3064 VDD.n1106 VDD.n1104 136.8
R3065 VDD.n1102 VDD.n1085 136.8
R3066 VDD.n1098 VDD.n1096 136.8
R3067 VDD.n1094 VDD.n1087 136.8
R3068 VDD.n1078 VDD.n1076 136.8
R3069 VDD.n1126 VDD.n1076 136.8
R3070 VDD.n1126 VDD.n1074 136.8
R3071 VDD.n1130 VDD.n1074 136.8
R3072 VDD.n1130 VDD.n1071 136.8
R3073 VDD.n1135 VDD.n1071 136.8
R3074 VDD.n1135 VDD.n1069 136.8
R3075 VDD.n1139 VDD.n1069 136.8
R3076 VDD.n1139 VDD.n1057 136.8
R3077 VDD.n1156 VDD.n1057 136.8
R3078 VDD.n1156 VDD.n1055 136.8
R3079 VDD.n1160 VDD.n1055 136.8
R3080 VDD.n1160 VDD.n1046 136.8
R3081 VDD.n1177 VDD.n1046 136.8
R3082 VDD.n1177 VDD.n1044 136.8
R3083 VDD.n1181 VDD.n1044 136.8
R3084 VDD.n1181 VDD.n1035 136.8
R3085 VDD.n1198 VDD.n1035 136.8
R3086 VDD.n1198 VDD.n1033 136.8
R3087 VDD.n1203 VDD.n1033 136.8
R3088 VDD.n1203 VDD.n1024 136.8
R3089 VDD.n1220 VDD.n1024 136.8
R3090 VDD.n1221 VDD.n1220 136.8
R3091 VDD.n1221 VDD.n1021 136.8
R3092 VDD.n1022 VDD.n1021 136.8
R3093 VDD.n1226 VDD.n1022 136.8
R3094 VDD.n1226 VDD.n978 136.8
R3095 VDD.n1244 VDD.n978 136.8
R3096 VDD.n1244 VDD.n975 136.8
R3097 VDD.n1008 VDD.n1007 136.8
R3098 VDD.n1004 VDD.n1003 136.8
R3099 VDD.n1000 VDD.n999 136.8
R3100 VDD.n996 VDD.n995 136.8
R3101 VDD.n992 VDD.n991 136.8
R3102 VDD.n988 VDD.n987 136.8
R3103 VDD.n984 VDD.n983 136.8
R3104 VDD.n1248 VDD.n974 136.8
R3105 VDD.n801 VDD.n799 136.8
R3106 VDD.n908 VDD.n907 136.8
R3107 VDD.n905 VDD.n284 136.8
R3108 VDD.n900 VDD.n899 136.8
R3109 VDD.n897 VDD.n288 136.8
R3110 VDD.n893 VDD.n892 136.8
R3111 VDD.n890 VDD.n291 136.8
R3112 VDD.n886 VDD.n885 136.8
R3113 VDD.n883 VDD.n294 136.8
R3114 VDD.n879 VDD.n878 136.8
R3115 VDD.n876 VDD.n297 136.8
R3116 VDD.n872 VDD.n871 136.8
R3117 VDD.n869 VDD.n300 136.8
R3118 VDD.n865 VDD.n864 136.8
R3119 VDD.n862 VDD.n303 136.8
R3120 VDD.n858 VDD.n857 136.8
R3121 VDD.n855 VDD.n306 136.8
R3122 VDD.n851 VDD.n850 136.8
R3123 VDD.n848 VDD.n309 136.8
R3124 VDD.n844 VDD.n843 136.8
R3125 VDD.n841 VDD.n312 136.8
R3126 VDD.n837 VDD.n836 136.8
R3127 VDD.n834 VDD.n315 136.8
R3128 VDD.n830 VDD.n829 136.8
R3129 VDD.n827 VDD.n318 136.8
R3130 VDD.n823 VDD.n822 136.8
R3131 VDD.n820 VDD.n321 136.8
R3132 VDD.n816 VDD.n815 136.8
R3133 VDD.n792 VDD.n326 136.8
R3134 VDD.n809 VDD.n326 136.8
R3135 VDD.n809 VDD.n324 136.8
R3136 VDD.n681 VDD.n680 136.8
R3137 VDD.n683 VDD.n681 136.8
R3138 VDD.n687 VDD.n676 136.8
R3139 VDD.n691 VDD.n689 136.8
R3140 VDD.n695 VDD.n674 136.8
R3141 VDD.n699 VDD.n697 136.8
R3142 VDD.n703 VDD.n672 136.8
R3143 VDD.n707 VDD.n705 136.8
R3144 VDD.n711 VDD.n670 136.8
R3145 VDD.n715 VDD.n713 136.8
R3146 VDD.n719 VDD.n668 136.8
R3147 VDD.n723 VDD.n721 136.8
R3148 VDD.n727 VDD.n666 136.8
R3149 VDD.n731 VDD.n729 136.8
R3150 VDD.n735 VDD.n664 136.8
R3151 VDD.n739 VDD.n737 136.8
R3152 VDD.n743 VDD.n662 136.8
R3153 VDD.n747 VDD.n745 136.8
R3154 VDD.n751 VDD.n660 136.8
R3155 VDD.n755 VDD.n753 136.8
R3156 VDD.n759 VDD.n658 136.8
R3157 VDD.n763 VDD.n761 136.8
R3158 VDD.n767 VDD.n656 136.8
R3159 VDD.n771 VDD.n769 136.8
R3160 VDD.n775 VDD.n654 136.8
R3161 VDD.n779 VDD.n777 136.8
R3162 VDD.n783 VDD.n652 136.8
R3163 VDD.n786 VDD.n785 136.8
R3164 VDD.n788 VDD.n649 136.8
R3165 VDD.n795 VDD.n328 136.8
R3166 VDD.n807 VDD.n328 136.8
R3167 VDD.n807 VDD.n329 136.8
R3168 VDD.n633 VDD.n632 136.8
R3169 VDD.n629 VDD.n628 136.8
R3170 VDD.n625 VDD.n624 136.8
R3171 VDD.n621 VDD.n620 136.8
R3172 VDD.n617 VDD.n616 136.8
R3173 VDD.n613 VDD.n612 136.8
R3174 VDD.n609 VDD.n608 136.8
R3175 VDD.n605 VDD.n604 136.8
R3176 VDD.n601 VDD.n600 136.8
R3177 VDD.n597 VDD.n596 136.8
R3178 VDD.n593 VDD.n592 136.8
R3179 VDD.n589 VDD.n588 136.8
R3180 VDD.n585 VDD.n584 136.8
R3181 VDD.n581 VDD.n580 136.8
R3182 VDD.n577 VDD.n576 136.8
R3183 VDD.n573 VDD.n572 136.8
R3184 VDD.n569 VDD.n568 136.8
R3185 VDD.n565 VDD.n564 136.8
R3186 VDD.n561 VDD.n560 136.8
R3187 VDD.n557 VDD.n556 136.8
R3188 VDD.n553 VDD.n552 136.8
R3189 VDD.n549 VDD.n548 136.8
R3190 VDD.n545 VDD.n544 136.8
R3191 VDD.n541 VDD.n540 136.8
R3192 VDD.n537 VDD.n536 136.8
R3193 VDD.n533 VDD.n532 136.8
R3194 VDD.n529 VDD.n528 136.8
R3195 VDD.n525 VDD.n361 136.8
R3196 VDD.n519 VDD.n365 136.8
R3197 VDD.n641 VDD.n365 136.8
R3198 VDD.n641 VDD.n362 136.8
R3199 VDD.n406 VDD.n405 136.8
R3200 VDD.n408 VDD.n406 136.8
R3201 VDD.n414 VDD.n399 136.8
R3202 VDD.n418 VDD.n416 136.8
R3203 VDD.n422 VDD.n396 136.8
R3204 VDD.n426 VDD.n424 136.8
R3205 VDD.n430 VDD.n394 136.8
R3206 VDD.n434 VDD.n432 136.8
R3207 VDD.n438 VDD.n392 136.8
R3208 VDD.n442 VDD.n440 136.8
R3209 VDD.n446 VDD.n390 136.8
R3210 VDD.n450 VDD.n448 136.8
R3211 VDD.n454 VDD.n388 136.8
R3212 VDD.n458 VDD.n456 136.8
R3213 VDD.n462 VDD.n386 136.8
R3214 VDD.n466 VDD.n464 136.8
R3215 VDD.n470 VDD.n384 136.8
R3216 VDD.n474 VDD.n472 136.8
R3217 VDD.n478 VDD.n382 136.8
R3218 VDD.n482 VDD.n480 136.8
R3219 VDD.n486 VDD.n380 136.8
R3220 VDD.n490 VDD.n488 136.8
R3221 VDD.n494 VDD.n378 136.8
R3222 VDD.n498 VDD.n496 136.8
R3223 VDD.n502 VDD.n376 136.8
R3224 VDD.n506 VDD.n504 136.8
R3225 VDD.n510 VDD.n374 136.8
R3226 VDD.n513 VDD.n512 136.8
R3227 VDD.n515 VDD.n371 136.8
R3228 VDD.n522 VDD.n366 136.8
R3229 VDD.n639 VDD.n366 136.8
R3230 VDD.n639 VDD.n367 136.8
R3231 VDD.n188 VDD.n187 136.8
R3232 VDD.n193 VDD.n190 136.8
R3233 VDD.n191 VDD.n46 136.8
R3234 VDD.n48 VDD.n47 136.8
R3235 VDD.n59 VDD.n52 136.8
R3236 VDD.n54 VDD.n53 136.8
R3237 VDD.n261 VDD.n57 136.8
R3238 VDD.n256 VDD.n68 136.8
R3239 VDD.n252 VDD.n68 136.8
R3240 VDD.n252 VDD.n203 136.8
R3241 VDD.n221 VDD.n219 136.8
R3242 VDD.n225 VDD.n214 136.8
R3243 VDD.n229 VDD.n227 136.8
R3244 VDD.n233 VDD.n212 136.8
R3245 VDD.n237 VDD.n235 136.8
R3246 VDD.n241 VDD.n210 136.8
R3247 VDD.n245 VDD.n243 136.8
R3248 VDD.n258 VDD.n64 136.8
R3249 VDD.n204 VDD.n64 136.8
R3250 VDD.n249 VDD.n204 136.8
R3251 VDD.n98 VDD.n97 136.8
R3252 VDD.n101 VDD.n100 136.8
R3253 VDD.n106 VDD.n103 136.8
R3254 VDD.n104 VDD.n74 136.8
R3255 VDD.n76 VDD.n75 136.8
R3256 VDD.n86 VDD.n79 136.8
R3257 VDD.n81 VDD.n80 136.8
R3258 VDD.n169 VDD.n93 136.8
R3259 VDD.n165 VDD.n93 136.8
R3260 VDD.n165 VDD.n117 136.8
R3261 VDD.n134 VDD.n132 136.8
R3262 VDD.n138 VDD.n127 136.8
R3263 VDD.n142 VDD.n140 136.8
R3264 VDD.n146 VDD.n125 136.8
R3265 VDD.n150 VDD.n148 136.8
R3266 VDD.n154 VDD.n123 136.8
R3267 VDD.n158 VDD.n156 136.8
R3268 VDD.n171 VDD.n84 136.8
R3269 VDD.n118 VDD.n84 136.8
R3270 VDD.n162 VDD.n118 136.8
R3271 VDD.n1403 VDD.t36 104.135
R3272 VDD.t19 VDD.n1411 104.135
R3273 VDD.n1396 VDD.t5 96.8274
R3274 VDD.t26 VDD.n1418 96.8274
R3275 VDD.t5 VDD.n1395 78.5582
R3276 VDD.n1419 VDD.t26 78.5582
R3277 VDD.n1373 VDD.t7 74.9043
R3278 VDD.t22 VDD.n1424 74.9043
R3279 VDD.n257 VDD.n63 73.592
R3280 VDD.n250 VDD.n205 73.592
R3281 VDD.n170 VDD.n90 73.592
R3282 VDD.n163 VDD.n119 73.592
R3283 VDD.n1406 VDD.t36 71.2505
R3284 VDD.n1412 VDD.t19 71.2505
R3285 VDD.n1425 VDD.n30 68.6629
R3286 VDD.n1371 VDD.n1370 68.6629
R3287 VDD.n1288 VDD.n1287 67.5326
R3288 VDD.n1288 VDD.n1250 67.5326
R3289 VDD.n1288 VDD.n1251 67.5326
R3290 VDD.n1288 VDD.n1252 67.5326
R3291 VDD.n1288 VDD.n1253 67.5326
R3292 VDD.n1288 VDD.n1254 67.5326
R3293 VDD.n1288 VDD.n1255 67.5326
R3294 VDD.n1289 VDD.n1288 67.5326
R3295 VDD.n1328 VDD.n954 67.5326
R3296 VDD.n1328 VDD.n955 67.5326
R3297 VDD.n1328 VDD.n956 67.5326
R3298 VDD.n1328 VDD.n957 67.5326
R3299 VDD.n1328 VDD.n958 67.5326
R3300 VDD.n1328 VDD.n959 67.5326
R3301 VDD.n1328 VDD.n960 67.5326
R3302 VDD.n1328 VDD.n1327 67.5326
R3303 VDD.n1249 VDD.n973 67.5326
R3304 VDD.n1249 VDD.n972 67.5326
R3305 VDD.n1249 VDD.n971 67.5326
R3306 VDD.n1249 VDD.n970 67.5326
R3307 VDD.n1249 VDD.n969 67.5326
R3308 VDD.n1249 VDD.n968 67.5326
R3309 VDD.n1249 VDD.n967 67.5326
R3310 VDD.n1249 VDD.n966 67.5326
R3311 VDD.n1079 VDD.n1077 67.5326
R3312 VDD.n1081 VDD.n1077 67.5326
R3313 VDD.n1111 VDD.n1077 67.5326
R3314 VDD.n1105 VDD.n1077 67.5326
R3315 VDD.n1103 VDD.n1077 67.5326
R3316 VDD.n1097 VDD.n1077 67.5326
R3317 VDD.n1095 VDD.n1077 67.5326
R3318 VDD.n1089 VDD.n1077 67.5326
R3319 VDD.n679 VDD.n648 67.5326
R3320 VDD.n682 VDD.n648 67.5326
R3321 VDD.n688 VDD.n648 67.5326
R3322 VDD.n690 VDD.n648 67.5326
R3323 VDD.n696 VDD.n648 67.5326
R3324 VDD.n698 VDD.n648 67.5326
R3325 VDD.n704 VDD.n648 67.5326
R3326 VDD.n706 VDD.n648 67.5326
R3327 VDD.n712 VDD.n648 67.5326
R3328 VDD.n714 VDD.n648 67.5326
R3329 VDD.n720 VDD.n648 67.5326
R3330 VDD.n722 VDD.n648 67.5326
R3331 VDD.n728 VDD.n648 67.5326
R3332 VDD.n730 VDD.n648 67.5326
R3333 VDD.n736 VDD.n648 67.5326
R3334 VDD.n738 VDD.n648 67.5326
R3335 VDD.n744 VDD.n648 67.5326
R3336 VDD.n746 VDD.n648 67.5326
R3337 VDD.n752 VDD.n648 67.5326
R3338 VDD.n754 VDD.n648 67.5326
R3339 VDD.n760 VDD.n648 67.5326
R3340 VDD.n762 VDD.n648 67.5326
R3341 VDD.n768 VDD.n648 67.5326
R3342 VDD.n770 VDD.n648 67.5326
R3343 VDD.n776 VDD.n648 67.5326
R3344 VDD.n778 VDD.n648 67.5326
R3345 VDD.n784 VDD.n648 67.5326
R3346 VDD.n787 VDD.n648 67.5326
R3347 VDD.n814 VDD.n283 67.5326
R3348 VDD.n323 VDD.n283 67.5326
R3349 VDD.n821 VDD.n283 67.5326
R3350 VDD.n320 VDD.n283 67.5326
R3351 VDD.n828 VDD.n283 67.5326
R3352 VDD.n317 VDD.n283 67.5326
R3353 VDD.n835 VDD.n283 67.5326
R3354 VDD.n314 VDD.n283 67.5326
R3355 VDD.n842 VDD.n283 67.5326
R3356 VDD.n311 VDD.n283 67.5326
R3357 VDD.n849 VDD.n283 67.5326
R3358 VDD.n308 VDD.n283 67.5326
R3359 VDD.n856 VDD.n283 67.5326
R3360 VDD.n305 VDD.n283 67.5326
R3361 VDD.n863 VDD.n283 67.5326
R3362 VDD.n302 VDD.n283 67.5326
R3363 VDD.n870 VDD.n283 67.5326
R3364 VDD.n299 VDD.n283 67.5326
R3365 VDD.n877 VDD.n283 67.5326
R3366 VDD.n296 VDD.n283 67.5326
R3367 VDD.n884 VDD.n283 67.5326
R3368 VDD.n293 VDD.n283 67.5326
R3369 VDD.n891 VDD.n283 67.5326
R3370 VDD.n290 VDD.n283 67.5326
R3371 VDD.n898 VDD.n283 67.5326
R3372 VDD.n287 VDD.n283 67.5326
R3373 VDD.n906 VDD.n283 67.5326
R3374 VDD.n283 VDD.n282 67.5326
R3375 VDD.n802 VDD.n283 67.5326
R3376 VDD.n647 VDD.n646 67.5326
R3377 VDD.n647 VDD.n360 67.5326
R3378 VDD.n647 VDD.n359 67.5326
R3379 VDD.n647 VDD.n358 67.5326
R3380 VDD.n647 VDD.n357 67.5326
R3381 VDD.n647 VDD.n356 67.5326
R3382 VDD.n647 VDD.n355 67.5326
R3383 VDD.n647 VDD.n354 67.5326
R3384 VDD.n647 VDD.n353 67.5326
R3385 VDD.n647 VDD.n352 67.5326
R3386 VDD.n647 VDD.n351 67.5326
R3387 VDD.n647 VDD.n350 67.5326
R3388 VDD.n647 VDD.n349 67.5326
R3389 VDD.n647 VDD.n348 67.5326
R3390 VDD.n647 VDD.n347 67.5326
R3391 VDD.n647 VDD.n346 67.5326
R3392 VDD.n647 VDD.n345 67.5326
R3393 VDD.n647 VDD.n344 67.5326
R3394 VDD.n647 VDD.n343 67.5326
R3395 VDD.n647 VDD.n342 67.5326
R3396 VDD.n647 VDD.n341 67.5326
R3397 VDD.n647 VDD.n340 67.5326
R3398 VDD.n647 VDD.n339 67.5326
R3399 VDD.n647 VDD.n338 67.5326
R3400 VDD.n647 VDD.n337 67.5326
R3401 VDD.n647 VDD.n336 67.5326
R3402 VDD.n647 VDD.n335 67.5326
R3403 VDD.n647 VDD.n334 67.5326
R3404 VDD.n647 VDD.n333 67.5326
R3405 VDD.n404 VDD.n370 67.5326
R3406 VDD.n407 VDD.n370 67.5326
R3407 VDD.n415 VDD.n370 67.5326
R3408 VDD.n417 VDD.n370 67.5326
R3409 VDD.n423 VDD.n370 67.5326
R3410 VDD.n425 VDD.n370 67.5326
R3411 VDD.n431 VDD.n370 67.5326
R3412 VDD.n433 VDD.n370 67.5326
R3413 VDD.n439 VDD.n370 67.5326
R3414 VDD.n441 VDD.n370 67.5326
R3415 VDD.n447 VDD.n370 67.5326
R3416 VDD.n449 VDD.n370 67.5326
R3417 VDD.n455 VDD.n370 67.5326
R3418 VDD.n457 VDD.n370 67.5326
R3419 VDD.n463 VDD.n370 67.5326
R3420 VDD.n465 VDD.n370 67.5326
R3421 VDD.n471 VDD.n370 67.5326
R3422 VDD.n473 VDD.n370 67.5326
R3423 VDD.n479 VDD.n370 67.5326
R3424 VDD.n481 VDD.n370 67.5326
R3425 VDD.n487 VDD.n370 67.5326
R3426 VDD.n489 VDD.n370 67.5326
R3427 VDD.n495 VDD.n370 67.5326
R3428 VDD.n497 VDD.n370 67.5326
R3429 VDD.n503 VDD.n370 67.5326
R3430 VDD.n505 VDD.n370 67.5326
R3431 VDD.n511 VDD.n370 67.5326
R3432 VDD.n514 VDD.n370 67.5326
R3433 VDD.n244 VDD.n205 67.5326
R3434 VDD.n242 VDD.n205 67.5326
R3435 VDD.n236 VDD.n205 67.5326
R3436 VDD.n234 VDD.n205 67.5326
R3437 VDD.n228 VDD.n205 67.5326
R3438 VDD.n226 VDD.n205 67.5326
R3439 VDD.n220 VDD.n205 67.5326
R3440 VDD.n218 VDD.n205 67.5326
R3441 VDD.n260 VDD.n63 67.5326
R3442 VDD.n63 VDD.n62 67.5326
R3443 VDD.n63 VDD.n61 67.5326
R3444 VDD.n63 VDD.n60 67.5326
R3445 VDD.n63 VDD.n58 67.5326
R3446 VDD.n192 VDD.n63 67.5326
R3447 VDD.n189 VDD.n63 67.5326
R3448 VDD.n186 VDD.n63 67.5326
R3449 VDD.n157 VDD.n119 67.5326
R3450 VDD.n155 VDD.n119 67.5326
R3451 VDD.n149 VDD.n119 67.5326
R3452 VDD.n147 VDD.n119 67.5326
R3453 VDD.n141 VDD.n119 67.5326
R3454 VDD.n139 VDD.n119 67.5326
R3455 VDD.n133 VDD.n119 67.5326
R3456 VDD.n131 VDD.n119 67.5326
R3457 VDD.n90 VDD.n89 67.5326
R3458 VDD.n90 VDD.n88 67.5326
R3459 VDD.n90 VDD.n87 67.5326
R3460 VDD.n90 VDD.n85 67.5326
R3461 VDD.n105 VDD.n90 67.5326
R3462 VDD.n102 VDD.n90 67.5326
R3463 VDD.n99 VDD.n90 67.5326
R3464 VDD.n96 VDD.n90 67.5326
R3465 VDD.n1123 VDD.n1077 67.5192
R3466 VDD.n1249 VDD.n965 67.5192
R3467 VDD.n1288 VDD.n947 67.5192
R3468 VDD.n1328 VDD.n951 67.5192
R3469 VDD.n184 VDD.t3 51.6977
R3470 VDD.n50 VDD.t18 51.6066
R3471 VDD.n648 VDD.n647 51.228
R3472 VDD.n1327 VDD.n1326 49.9379
R3473 VDD.n1322 VDD.n960 49.9379
R3474 VDD.n1318 VDD.n959 49.9379
R3475 VDD.n1314 VDD.n958 49.9379
R3476 VDD.n1310 VDD.n957 49.9379
R3477 VDD.n1306 VDD.n956 49.9379
R3478 VDD.n1302 VDD.n955 49.9379
R3479 VDD.n1298 VDD.n954 49.9379
R3480 VDD.n1287 VDD.n1286 49.9379
R3481 VDD.n1281 VDD.n1250 49.9379
R3482 VDD.n1278 VDD.n1251 49.9379
R3483 VDD.n1274 VDD.n1252 49.9379
R3484 VDD.n1270 VDD.n1253 49.9379
R3485 VDD.n1266 VDD.n1254 49.9379
R3486 VDD.n1262 VDD.n1255 49.9379
R3487 VDD.n1289 VDD.n964 49.9379
R3488 VDD.n1287 VDD.n1257 49.9379
R3489 VDD.n1279 VDD.n1250 49.9379
R3490 VDD.n1275 VDD.n1251 49.9379
R3491 VDD.n1271 VDD.n1252 49.9379
R3492 VDD.n1267 VDD.n1253 49.9379
R3493 VDD.n1263 VDD.n1254 49.9379
R3494 VDD.n1259 VDD.n1255 49.9379
R3495 VDD.n1290 VDD.n1289 49.9379
R3496 VDD.n1301 VDD.n954 49.9379
R3497 VDD.n1305 VDD.n955 49.9379
R3498 VDD.n1309 VDD.n956 49.9379
R3499 VDD.n1313 VDD.n957 49.9379
R3500 VDD.n1317 VDD.n958 49.9379
R3501 VDD.n1321 VDD.n959 49.9379
R3502 VDD.n961 VDD.n960 49.9379
R3503 VDD.n1327 VDD.n952 49.9379
R3504 VDD.n1121 VDD.n1079 49.9379
R3505 VDD.n1116 VDD.n1081 49.9379
R3506 VDD.n1112 VDD.n1111 49.9379
R3507 VDD.n1105 VDD.n1083 49.9379
R3508 VDD.n1104 VDD.n1103 49.9379
R3509 VDD.n1097 VDD.n1085 49.9379
R3510 VDD.n1096 VDD.n1095 49.9379
R3511 VDD.n1089 VDD.n1087 49.9379
R3512 VDD.n981 VDD.n966 49.9379
R3513 VDD.n1007 VDD.n967 49.9379
R3514 VDD.n1003 VDD.n968 49.9379
R3515 VDD.n999 VDD.n969 49.9379
R3516 VDD.n995 VDD.n970 49.9379
R3517 VDD.n991 VDD.n971 49.9379
R3518 VDD.n987 VDD.n972 49.9379
R3519 VDD.n983 VDD.n973 49.9379
R3520 VDD.n974 VDD.n973 49.9379
R3521 VDD.n984 VDD.n972 49.9379
R3522 VDD.n988 VDD.n971 49.9379
R3523 VDD.n992 VDD.n970 49.9379
R3524 VDD.n996 VDD.n969 49.9379
R3525 VDD.n1000 VDD.n968 49.9379
R3526 VDD.n1004 VDD.n967 49.9379
R3527 VDD.n1008 VDD.n966 49.9379
R3528 VDD.n1118 VDD.n1079 49.9379
R3529 VDD.n1113 VDD.n1081 49.9379
R3530 VDD.n1111 VDD.n1110 49.9379
R3531 VDD.n1106 VDD.n1105 49.9379
R3532 VDD.n1103 VDD.n1102 49.9379
R3533 VDD.n1098 VDD.n1097 49.9379
R3534 VDD.n1095 VDD.n1094 49.9379
R3535 VDD.n1090 VDD.n1089 49.9379
R3536 VDD.n802 VDD.n801 49.9379
R3537 VDD.n908 VDD.n282 49.9379
R3538 VDD.n906 VDD.n905 49.9379
R3539 VDD.n900 VDD.n287 49.9379
R3540 VDD.n898 VDD.n897 49.9379
R3541 VDD.n893 VDD.n290 49.9379
R3542 VDD.n891 VDD.n890 49.9379
R3543 VDD.n886 VDD.n293 49.9379
R3544 VDD.n884 VDD.n883 49.9379
R3545 VDD.n879 VDD.n296 49.9379
R3546 VDD.n877 VDD.n876 49.9379
R3547 VDD.n872 VDD.n299 49.9379
R3548 VDD.n870 VDD.n869 49.9379
R3549 VDD.n865 VDD.n302 49.9379
R3550 VDD.n863 VDD.n862 49.9379
R3551 VDD.n858 VDD.n305 49.9379
R3552 VDD.n856 VDD.n855 49.9379
R3553 VDD.n851 VDD.n308 49.9379
R3554 VDD.n849 VDD.n848 49.9379
R3555 VDD.n844 VDD.n311 49.9379
R3556 VDD.n842 VDD.n841 49.9379
R3557 VDD.n837 VDD.n314 49.9379
R3558 VDD.n835 VDD.n834 49.9379
R3559 VDD.n830 VDD.n317 49.9379
R3560 VDD.n828 VDD.n827 49.9379
R3561 VDD.n823 VDD.n320 49.9379
R3562 VDD.n821 VDD.n820 49.9379
R3563 VDD.n816 VDD.n323 49.9379
R3564 VDD.n814 VDD.n813 49.9379
R3565 VDD.n679 VDD.n331 49.9379
R3566 VDD.n683 VDD.n682 49.9379
R3567 VDD.n688 VDD.n687 49.9379
R3568 VDD.n691 VDD.n690 49.9379
R3569 VDD.n696 VDD.n695 49.9379
R3570 VDD.n699 VDD.n698 49.9379
R3571 VDD.n704 VDD.n703 49.9379
R3572 VDD.n707 VDD.n706 49.9379
R3573 VDD.n712 VDD.n711 49.9379
R3574 VDD.n715 VDD.n714 49.9379
R3575 VDD.n720 VDD.n719 49.9379
R3576 VDD.n723 VDD.n722 49.9379
R3577 VDD.n728 VDD.n727 49.9379
R3578 VDD.n731 VDD.n730 49.9379
R3579 VDD.n736 VDD.n735 49.9379
R3580 VDD.n739 VDD.n738 49.9379
R3581 VDD.n744 VDD.n743 49.9379
R3582 VDD.n747 VDD.n746 49.9379
R3583 VDD.n752 VDD.n751 49.9379
R3584 VDD.n755 VDD.n754 49.9379
R3585 VDD.n760 VDD.n759 49.9379
R3586 VDD.n763 VDD.n762 49.9379
R3587 VDD.n768 VDD.n767 49.9379
R3588 VDD.n771 VDD.n770 49.9379
R3589 VDD.n776 VDD.n775 49.9379
R3590 VDD.n779 VDD.n778 49.9379
R3591 VDD.n784 VDD.n783 49.9379
R3592 VDD.n787 VDD.n786 49.9379
R3593 VDD.n680 VDD.n679 49.9379
R3594 VDD.n682 VDD.n676 49.9379
R3595 VDD.n689 VDD.n688 49.9379
R3596 VDD.n690 VDD.n674 49.9379
R3597 VDD.n697 VDD.n696 49.9379
R3598 VDD.n698 VDD.n672 49.9379
R3599 VDD.n705 VDD.n704 49.9379
R3600 VDD.n706 VDD.n670 49.9379
R3601 VDD.n713 VDD.n712 49.9379
R3602 VDD.n714 VDD.n668 49.9379
R3603 VDD.n721 VDD.n720 49.9379
R3604 VDD.n722 VDD.n666 49.9379
R3605 VDD.n729 VDD.n728 49.9379
R3606 VDD.n730 VDD.n664 49.9379
R3607 VDD.n737 VDD.n736 49.9379
R3608 VDD.n738 VDD.n662 49.9379
R3609 VDD.n745 VDD.n744 49.9379
R3610 VDD.n746 VDD.n660 49.9379
R3611 VDD.n753 VDD.n752 49.9379
R3612 VDD.n754 VDD.n658 49.9379
R3613 VDD.n761 VDD.n760 49.9379
R3614 VDD.n762 VDD.n656 49.9379
R3615 VDD.n769 VDD.n768 49.9379
R3616 VDD.n770 VDD.n654 49.9379
R3617 VDD.n777 VDD.n776 49.9379
R3618 VDD.n778 VDD.n652 49.9379
R3619 VDD.n785 VDD.n784 49.9379
R3620 VDD.n788 VDD.n787 49.9379
R3621 VDD.n815 VDD.n814 49.9379
R3622 VDD.n323 VDD.n321 49.9379
R3623 VDD.n822 VDD.n821 49.9379
R3624 VDD.n320 VDD.n318 49.9379
R3625 VDD.n829 VDD.n828 49.9379
R3626 VDD.n317 VDD.n315 49.9379
R3627 VDD.n836 VDD.n835 49.9379
R3628 VDD.n314 VDD.n312 49.9379
R3629 VDD.n843 VDD.n842 49.9379
R3630 VDD.n311 VDD.n309 49.9379
R3631 VDD.n850 VDD.n849 49.9379
R3632 VDD.n308 VDD.n306 49.9379
R3633 VDD.n857 VDD.n856 49.9379
R3634 VDD.n305 VDD.n303 49.9379
R3635 VDD.n864 VDD.n863 49.9379
R3636 VDD.n302 VDD.n300 49.9379
R3637 VDD.n871 VDD.n870 49.9379
R3638 VDD.n299 VDD.n297 49.9379
R3639 VDD.n878 VDD.n877 49.9379
R3640 VDD.n296 VDD.n294 49.9379
R3641 VDD.n885 VDD.n884 49.9379
R3642 VDD.n293 VDD.n291 49.9379
R3643 VDD.n892 VDD.n891 49.9379
R3644 VDD.n290 VDD.n288 49.9379
R3645 VDD.n899 VDD.n898 49.9379
R3646 VDD.n287 VDD.n284 49.9379
R3647 VDD.n907 VDD.n906 49.9379
R3648 VDD.n799 VDD.n282 49.9379
R3649 VDD.n803 VDD.n802 49.9379
R3650 VDD.n633 VDD.n333 49.9379
R3651 VDD.n629 VDD.n334 49.9379
R3652 VDD.n625 VDD.n335 49.9379
R3653 VDD.n621 VDD.n336 49.9379
R3654 VDD.n617 VDD.n337 49.9379
R3655 VDD.n613 VDD.n338 49.9379
R3656 VDD.n609 VDD.n339 49.9379
R3657 VDD.n605 VDD.n340 49.9379
R3658 VDD.n601 VDD.n341 49.9379
R3659 VDD.n597 VDD.n342 49.9379
R3660 VDD.n593 VDD.n343 49.9379
R3661 VDD.n589 VDD.n344 49.9379
R3662 VDD.n585 VDD.n345 49.9379
R3663 VDD.n581 VDD.n346 49.9379
R3664 VDD.n577 VDD.n347 49.9379
R3665 VDD.n573 VDD.n348 49.9379
R3666 VDD.n569 VDD.n349 49.9379
R3667 VDD.n565 VDD.n350 49.9379
R3668 VDD.n561 VDD.n351 49.9379
R3669 VDD.n557 VDD.n352 49.9379
R3670 VDD.n553 VDD.n353 49.9379
R3671 VDD.n549 VDD.n354 49.9379
R3672 VDD.n545 VDD.n355 49.9379
R3673 VDD.n541 VDD.n356 49.9379
R3674 VDD.n537 VDD.n357 49.9379
R3675 VDD.n533 VDD.n358 49.9379
R3676 VDD.n529 VDD.n359 49.9379
R3677 VDD.n525 VDD.n360 49.9379
R3678 VDD.n646 VDD.n645 49.9379
R3679 VDD.n404 VDD.n369 49.9379
R3680 VDD.n408 VDD.n407 49.9379
R3681 VDD.n415 VDD.n414 49.9379
R3682 VDD.n418 VDD.n417 49.9379
R3683 VDD.n423 VDD.n422 49.9379
R3684 VDD.n426 VDD.n425 49.9379
R3685 VDD.n431 VDD.n430 49.9379
R3686 VDD.n434 VDD.n433 49.9379
R3687 VDD.n439 VDD.n438 49.9379
R3688 VDD.n442 VDD.n441 49.9379
R3689 VDD.n447 VDD.n446 49.9379
R3690 VDD.n450 VDD.n449 49.9379
R3691 VDD.n455 VDD.n454 49.9379
R3692 VDD.n458 VDD.n457 49.9379
R3693 VDD.n463 VDD.n462 49.9379
R3694 VDD.n466 VDD.n465 49.9379
R3695 VDD.n471 VDD.n470 49.9379
R3696 VDD.n474 VDD.n473 49.9379
R3697 VDD.n479 VDD.n478 49.9379
R3698 VDD.n482 VDD.n481 49.9379
R3699 VDD.n487 VDD.n486 49.9379
R3700 VDD.n490 VDD.n489 49.9379
R3701 VDD.n495 VDD.n494 49.9379
R3702 VDD.n498 VDD.n497 49.9379
R3703 VDD.n503 VDD.n502 49.9379
R3704 VDD.n506 VDD.n505 49.9379
R3705 VDD.n511 VDD.n510 49.9379
R3706 VDD.n514 VDD.n513 49.9379
R3707 VDD.n646 VDD.n361 49.9379
R3708 VDD.n528 VDD.n360 49.9379
R3709 VDD.n532 VDD.n359 49.9379
R3710 VDD.n536 VDD.n358 49.9379
R3711 VDD.n540 VDD.n357 49.9379
R3712 VDD.n544 VDD.n356 49.9379
R3713 VDD.n548 VDD.n355 49.9379
R3714 VDD.n552 VDD.n354 49.9379
R3715 VDD.n556 VDD.n353 49.9379
R3716 VDD.n560 VDD.n352 49.9379
R3717 VDD.n564 VDD.n351 49.9379
R3718 VDD.n568 VDD.n350 49.9379
R3719 VDD.n572 VDD.n349 49.9379
R3720 VDD.n576 VDD.n348 49.9379
R3721 VDD.n580 VDD.n347 49.9379
R3722 VDD.n584 VDD.n346 49.9379
R3723 VDD.n588 VDD.n345 49.9379
R3724 VDD.n592 VDD.n344 49.9379
R3725 VDD.n596 VDD.n343 49.9379
R3726 VDD.n600 VDD.n342 49.9379
R3727 VDD.n604 VDD.n341 49.9379
R3728 VDD.n608 VDD.n340 49.9379
R3729 VDD.n612 VDD.n339 49.9379
R3730 VDD.n616 VDD.n338 49.9379
R3731 VDD.n620 VDD.n337 49.9379
R3732 VDD.n624 VDD.n336 49.9379
R3733 VDD.n628 VDD.n335 49.9379
R3734 VDD.n632 VDD.n334 49.9379
R3735 VDD.n635 VDD.n333 49.9379
R3736 VDD.n405 VDD.n404 49.9379
R3737 VDD.n407 VDD.n399 49.9379
R3738 VDD.n416 VDD.n415 49.9379
R3739 VDD.n417 VDD.n396 49.9379
R3740 VDD.n424 VDD.n423 49.9379
R3741 VDD.n425 VDD.n394 49.9379
R3742 VDD.n432 VDD.n431 49.9379
R3743 VDD.n433 VDD.n392 49.9379
R3744 VDD.n440 VDD.n439 49.9379
R3745 VDD.n441 VDD.n390 49.9379
R3746 VDD.n448 VDD.n447 49.9379
R3747 VDD.n449 VDD.n388 49.9379
R3748 VDD.n456 VDD.n455 49.9379
R3749 VDD.n457 VDD.n386 49.9379
R3750 VDD.n464 VDD.n463 49.9379
R3751 VDD.n465 VDD.n384 49.9379
R3752 VDD.n472 VDD.n471 49.9379
R3753 VDD.n473 VDD.n382 49.9379
R3754 VDD.n480 VDD.n479 49.9379
R3755 VDD.n481 VDD.n380 49.9379
R3756 VDD.n488 VDD.n487 49.9379
R3757 VDD.n489 VDD.n378 49.9379
R3758 VDD.n496 VDD.n495 49.9379
R3759 VDD.n497 VDD.n376 49.9379
R3760 VDD.n504 VDD.n503 49.9379
R3761 VDD.n505 VDD.n374 49.9379
R3762 VDD.n512 VDD.n511 49.9379
R3763 VDD.n515 VDD.n514 49.9379
R3764 VDD.n187 VDD.n186 49.9379
R3765 VDD.n190 VDD.n189 49.9379
R3766 VDD.n192 VDD.n191 49.9379
R3767 VDD.n58 VDD.n47 49.9379
R3768 VDD.n60 VDD.n59 49.9379
R3769 VDD.n61 VDD.n53 49.9379
R3770 VDD.n62 VDD.n57 49.9379
R3771 VDD.n260 VDD.n259 49.9379
R3772 VDD.n219 VDD.n218 49.9379
R3773 VDD.n220 VDD.n214 49.9379
R3774 VDD.n227 VDD.n226 49.9379
R3775 VDD.n228 VDD.n212 49.9379
R3776 VDD.n235 VDD.n234 49.9379
R3777 VDD.n236 VDD.n210 49.9379
R3778 VDD.n243 VDD.n242 49.9379
R3779 VDD.n244 VDD.n206 49.9379
R3780 VDD.n245 VDD.n244 49.9379
R3781 VDD.n242 VDD.n241 49.9379
R3782 VDD.n237 VDD.n236 49.9379
R3783 VDD.n234 VDD.n233 49.9379
R3784 VDD.n229 VDD.n228 49.9379
R3785 VDD.n226 VDD.n225 49.9379
R3786 VDD.n221 VDD.n220 49.9379
R3787 VDD.n218 VDD.n217 49.9379
R3788 VDD.n261 VDD.n260 49.9379
R3789 VDD.n62 VDD.n54 49.9379
R3790 VDD.n61 VDD.n52 49.9379
R3791 VDD.n60 VDD.n48 49.9379
R3792 VDD.n58 VDD.n46 49.9379
R3793 VDD.n193 VDD.n192 49.9379
R3794 VDD.n189 VDD.n188 49.9379
R3795 VDD.n186 VDD.n67 49.9379
R3796 VDD.n97 VDD.n96 49.9379
R3797 VDD.n100 VDD.n99 49.9379
R3798 VDD.n103 VDD.n102 49.9379
R3799 VDD.n105 VDD.n104 49.9379
R3800 VDD.n85 VDD.n75 49.9379
R3801 VDD.n87 VDD.n86 49.9379
R3802 VDD.n88 VDD.n80 49.9379
R3803 VDD.n89 VDD.n82 49.9379
R3804 VDD.n132 VDD.n131 49.9379
R3805 VDD.n133 VDD.n127 49.9379
R3806 VDD.n140 VDD.n139 49.9379
R3807 VDD.n141 VDD.n125 49.9379
R3808 VDD.n148 VDD.n147 49.9379
R3809 VDD.n149 VDD.n123 49.9379
R3810 VDD.n156 VDD.n155 49.9379
R3811 VDD.n157 VDD.n120 49.9379
R3812 VDD.n158 VDD.n157 49.9379
R3813 VDD.n155 VDD.n154 49.9379
R3814 VDD.n150 VDD.n149 49.9379
R3815 VDD.n147 VDD.n146 49.9379
R3816 VDD.n142 VDD.n141 49.9379
R3817 VDD.n139 VDD.n138 49.9379
R3818 VDD.n134 VDD.n133 49.9379
R3819 VDD.n131 VDD.n130 49.9379
R3820 VDD.n89 VDD.n81 49.9379
R3821 VDD.n88 VDD.n79 49.9379
R3822 VDD.n87 VDD.n76 49.9379
R3823 VDD.n85 VDD.n74 49.9379
R3824 VDD.n106 VDD.n105 49.9379
R3825 VDD.n102 VDD.n101 49.9379
R3826 VDD.n99 VDD.n98 49.9379
R3827 VDD.n96 VDD.n92 49.9379
R3828 VDD.n65 VDD.n56 44.5872
R3829 VDD.n248 VDD.n247 44.5872
R3830 VDD.n216 VDD.n202 44.5872
R3831 VDD.n255 VDD.n201 44.5872
R3832 VDD.n173 VDD.n172 44.5872
R3833 VDD.n161 VDD.n160 44.5872
R3834 VDD.n129 VDD.n116 44.5872
R3835 VDD.n168 VDD.n115 44.5872
R3836 VDD.n257 VDD.n66 43.7905
R3837 VDD.n251 VDD.n250 43.7905
R3838 VDD.n170 VDD.n91 43.7905
R3839 VDD.n164 VDD.n163 43.7905
R3840 VDD.n1124 VDD.n1123 42.6439
R3841 VDD.n1125 VDD.n1124 42.6439
R3842 VDD.n1125 VDD.n1073 42.6439
R3843 VDD.n1131 VDD.n1073 42.6439
R3844 VDD.n1132 VDD.n1131 42.6439
R3845 VDD.n1134 VDD.n1132 42.6439
R3846 VDD.n1134 VDD.n1068 42.6439
R3847 VDD.n1140 VDD.n1068 42.6439
R3848 VDD.n1140 VDD.n1058 42.6439
R3849 VDD.n1155 VDD.n1058 42.6439
R3850 VDD.n1155 VDD.n1054 42.6439
R3851 VDD.n1161 VDD.n1054 42.6439
R3852 VDD.n1161 VDD.n1047 42.6439
R3853 VDD.n1176 VDD.n1047 42.6439
R3854 VDD.n1182 VDD.n1043 42.6439
R3855 VDD.n1182 VDD.n1036 42.6439
R3856 VDD.n1197 VDD.n1036 42.6439
R3857 VDD.n1197 VDD.n1032 42.6439
R3858 VDD.n1204 VDD.n1032 42.6439
R3859 VDD.n1204 VDD.n1025 42.6439
R3860 VDD.n1219 VDD.n1025 42.6439
R3861 VDD.n1219 VDD.n1020 42.6439
R3862 VDD.n1229 VDD.n1020 42.6439
R3863 VDD.n1229 VDD.n1228 42.6439
R3864 VDD.n1228 VDD.n1227 42.6439
R3865 VDD.n1227 VDD.n979 42.6439
R3866 VDD.n1243 VDD.n979 42.6439
R3867 VDD.n1243 VDD.n965 42.6439
R3868 VDD.n1335 VDD.n947 42.6439
R3869 VDD.n1335 VDD.n1334 42.6439
R3870 VDD.n1333 VDD.n951 42.6439
R3871 VDD.n805 VDD.n804 42.0272
R3872 VDD.n812 VDD.n811 42.0272
R3873 VDD.n791 VDD.n790 42.0272
R3874 VDD.n796 VDD.n330 42.0272
R3875 VDD.n523 VDD.n368 42.0272
R3876 VDD.n637 VDD.n636 42.0272
R3877 VDD.n644 VDD.n643 42.0272
R3878 VDD.n518 VDD.n517 42.0272
R3879 VDD.t15 VDD.n1043 41.4594
R3880 VDD.n1285 VDD.n943 39.8938
R3881 VDD.n953 VDD.n941 39.8938
R3882 VDD.n1299 VDD.n1296 39.8938
R3883 VDD.n1292 VDD.n963 39.8938
R3884 VDD.n1011 VDD.n1010 39.8938
R3885 VDD.n1247 VDD.n1246 39.8938
R3886 VDD.n1091 VDD.n1088 39.8938
R3887 VDD.n1120 VDD.n913 39.8938
R3888 VDD.n1369 VDD.n41 36.1417
R3889 VDD.n41 VDD.n39 36.1417
R3890 VDD.n1378 VDD.n39 36.1417
R3891 VDD.n1378 VDD.n1377 36.1417
R3892 VDD.n1377 VDD.n35 36.1417
R3893 VDD.n1393 VDD.n35 36.1417
R3894 VDD.n1393 VDD.n36 36.1417
R3895 VDD.n36 VDD.n32 36.1417
R3896 VDD.n32 VDD.n2 36.1417
R3897 VDD.n1471 VDD.n2 36.1417
R3898 VDD.n1471 VDD.n1470 36.1417
R3899 VDD.n1470 VDD.n5 36.1417
R3900 VDD.n8 VDD.n5 36.1417
R3901 VDD.n1463 VDD.n8 36.1417
R3902 VDD.n1463 VDD.n1462 36.1417
R3903 VDD.n1462 VDD.n11 36.1417
R3904 VDD.n1457 VDD.n11 36.1417
R3905 VDD.n1457 VDD.n1456 36.1417
R3906 VDD.n1456 VDD.n15 36.1417
R3907 VDD.n1450 VDD.n15 36.1417
R3908 VDD.n1450 VDD.n1449 36.1417
R3909 VDD.n1449 VDD.n20 36.1417
R3910 VDD.n1442 VDD.n20 36.1417
R3911 VDD.n1442 VDD.n1441 36.1417
R3912 VDD.n1441 VDD.n1440 36.1417
R3913 VDD.n1440 VDD.n26 36.1417
R3914 VDD.n1433 VDD.n26 36.1417
R3915 VDD.n1433 VDD.n1432 36.1417
R3916 VDD.n1432 VDD.n1426 36.1417
R3917 VDD.t11 VDD.n1374 34.712
R3918 VDD.n1423 VDD.t24 34.712
R3919 VDD.t9 VDD.n33 31.0582
R3920 VDD.t28 VDD.n1420 31.0582
R3921 VDD.n1353 VDD.n1352 27.1064
R3922 VDD.n1345 VDD.n926 27.1064
R3923 VDD.n1062 VDD.n927 27.1064
R3924 VDD.n1146 VDD.n1145 27.1064
R3925 VDD.n1150 VDD.n1149 27.1064
R3926 VDD.n1167 VDD.n1166 27.1064
R3927 VDD.n1171 VDD.n1170 27.1064
R3928 VDD.n1188 VDD.n1187 27.1064
R3929 VDD.n1192 VDD.n1191 27.1064
R3930 VDD.n1210 VDD.n1209 27.1064
R3931 VDD.n1214 VDD.n1213 27.1064
R3932 VDD.n1235 VDD.n1234 27.1064
R3933 VDD.n1342 VDD.n938 27.1064
R3934 VDD.n521 VDD.n370 25.1978
R3935 VDD.n647 VDD.n332 25.1978
R3936 VDD.n794 VDD.n648 25.1978
R3937 VDD.n327 VDD.n283 25.1978
R3938 VDD.n919 VDD.n914 22.5471
R3939 VDD.t13 VDD.n1333 22.5067
R3940 VDD.t17 VDD.n66 21.8955
R3941 VDD.n251 VDD.t17 21.8955
R3942 VDD.t2 VDD.n91 21.8955
R3943 VDD.n164 VDD.t2 21.8955
R3944 VDD.n1334 VDD.t13 20.1377
R3945 VDD.n1387 VDD.t6 17.8272
R3946 VDD.n1387 VDD.t31 17.8272
R3947 VDD.n1436 VDD.t29 17.8272
R3948 VDD.n1436 VDD.t25 17.8272
R3949 VDD.n1381 VDD.t12 17.8272
R3950 VDD.n1381 VDD.t10 17.8272
R3951 VDD.n1445 VDD.t35 17.8272
R3952 VDD.n1445 VDD.t27 17.8272
R3953 VDD.n1337 VDD.n944 15.3605
R3954 VDD.n1331 VDD.n941 15.3605
R3955 VDD.n962 VDD.n953 15.3605
R3956 VDD.n1325 VDD.n962 15.3605
R3957 VDD.n1325 VDD.n1324 15.3605
R3958 VDD.n1324 VDD.n1323 15.3605
R3959 VDD.n1323 VDD.n1320 15.3605
R3960 VDD.n1320 VDD.n1319 15.3605
R3961 VDD.n1319 VDD.n1316 15.3605
R3962 VDD.n1316 VDD.n1315 15.3605
R3963 VDD.n1315 VDD.n1312 15.3605
R3964 VDD.n1312 VDD.n1311 15.3605
R3965 VDD.n1311 VDD.n1308 15.3605
R3966 VDD.n1308 VDD.n1307 15.3605
R3967 VDD.n1307 VDD.n1304 15.3605
R3968 VDD.n1304 VDD.n1303 15.3605
R3969 VDD.n1303 VDD.n1300 15.3605
R3970 VDD.n1300 VDD.n1299 15.3605
R3971 VDD.n1293 VDD.n1292 15.3605
R3972 VDD.n1294 VDD.n1293 15.3605
R3973 VDD.n1295 VDD.n1294 15.3605
R3974 VDD.n1296 VDD.n1295 15.3605
R3975 VDD.n1285 VDD.n1284 15.3605
R3976 VDD.n1284 VDD.n1283 15.3605
R3977 VDD.n1283 VDD.n1282 15.3605
R3978 VDD.n1282 VDD.n1280 15.3605
R3979 VDD.n1280 VDD.n1277 15.3605
R3980 VDD.n1277 VDD.n1276 15.3605
R3981 VDD.n1276 VDD.n1273 15.3605
R3982 VDD.n1273 VDD.n1272 15.3605
R3983 VDD.n1272 VDD.n1269 15.3605
R3984 VDD.n1269 VDD.n1268 15.3605
R3985 VDD.n1268 VDD.n1265 15.3605
R3986 VDD.n1265 VDD.n1264 15.3605
R3987 VDD.n1264 VDD.n1261 15.3605
R3988 VDD.n1261 VDD.n1260 15.3605
R3989 VDD.n1260 VDD.n1258 15.3605
R3990 VDD.n1258 VDD.n963 15.3605
R3991 VDD.n1010 VDD.n1009 15.3605
R3992 VDD.n1009 VDD.n1006 15.3605
R3993 VDD.n1006 VDD.n1005 15.3605
R3994 VDD.n1005 VDD.n1002 15.3605
R3995 VDD.n1002 VDD.n1001 15.3605
R3996 VDD.n1001 VDD.n998 15.3605
R3997 VDD.n998 VDD.n997 15.3605
R3998 VDD.n997 VDD.n994 15.3605
R3999 VDD.n994 VDD.n993 15.3605
R4000 VDD.n993 VDD.n990 15.3605
R4001 VDD.n990 VDD.n989 15.3605
R4002 VDD.n989 VDD.n986 15.3605
R4003 VDD.n986 VDD.n985 15.3605
R4004 VDD.n985 VDD.n982 15.3605
R4005 VDD.n982 VDD.n976 15.3605
R4006 VDD.n1247 VDD.n976 15.3605
R4007 VDD.n1088 VDD.n1075 15.3605
R4008 VDD.n1127 VDD.n1075 15.3605
R4009 VDD.n1128 VDD.n1127 15.3605
R4010 VDD.n1129 VDD.n1128 15.3605
R4011 VDD.n1129 VDD.n1070 15.3605
R4012 VDD.n1136 VDD.n1070 15.3605
R4013 VDD.n1137 VDD.n1136 15.3605
R4014 VDD.n1138 VDD.n1137 15.3605
R4015 VDD.n1138 VDD.n1056 15.3605
R4016 VDD.n1157 VDD.n1056 15.3605
R4017 VDD.n1158 VDD.n1157 15.3605
R4018 VDD.n1159 VDD.n1158 15.3605
R4019 VDD.n1159 VDD.n1045 15.3605
R4020 VDD.n1178 VDD.n1045 15.3605
R4021 VDD.n1179 VDD.n1178 15.3605
R4022 VDD.n1180 VDD.n1179 15.3605
R4023 VDD.n1180 VDD.n1034 15.3605
R4024 VDD.n1199 VDD.n1034 15.3605
R4025 VDD.n1200 VDD.n1199 15.3605
R4026 VDD.n1202 VDD.n1200 15.3605
R4027 VDD.n1202 VDD.n1201 15.3605
R4028 VDD.n1201 VDD.n1023 15.3605
R4029 VDD.n1222 VDD.n1023 15.3605
R4030 VDD.n1223 VDD.n1222 15.3605
R4031 VDD.n1224 VDD.n1223 15.3605
R4032 VDD.n1225 VDD.n1224 15.3605
R4033 VDD.n1225 VDD.n977 15.3605
R4034 VDD.n1245 VDD.n977 15.3605
R4035 VDD.n1246 VDD.n1245 15.3605
R4036 VDD.n1120 VDD.n1119 15.3605
R4037 VDD.n1119 VDD.n1080 15.3605
R4038 VDD.n1115 VDD.n1080 15.3605
R4039 VDD.n1115 VDD.n1114 15.3605
R4040 VDD.n1114 VDD.n1082 15.3605
R4041 VDD.n1109 VDD.n1082 15.3605
R4042 VDD.n1109 VDD.n1108 15.3605
R4043 VDD.n1108 VDD.n1107 15.3605
R4044 VDD.n1107 VDD.n1084 15.3605
R4045 VDD.n1101 VDD.n1084 15.3605
R4046 VDD.n1101 VDD.n1100 15.3605
R4047 VDD.n1100 VDD.n1099 15.3605
R4048 VDD.n1099 VDD.n1086 15.3605
R4049 VDD.n1093 VDD.n1086 15.3605
R4050 VDD.n1093 VDD.n1092 15.3605
R4051 VDD.n1092 VDD.n1091 15.3605
R4052 VDD.n1357 VDD.n913 15.3605
R4053 VDD.n1357 VDD.n1356 15.3605
R4054 VDD.n1356 VDD.n917 15.3605
R4055 VDD.n1349 VDD.n917 15.3605
R4056 VDD.n1349 VDD.n1348 15.3605
R4057 VDD.n1348 VDD.n924 15.3605
R4058 VDD.n1066 VDD.n924 15.3605
R4059 VDD.n1142 VDD.n1066 15.3605
R4060 VDD.n1142 VDD.n1060 15.3605
R4061 VDD.n1153 VDD.n1060 15.3605
R4062 VDD.n1153 VDD.n1052 15.3605
R4063 VDD.n1163 VDD.n1052 15.3605
R4064 VDD.n1163 VDD.n1049 15.3605
R4065 VDD.n1174 VDD.n1049 15.3605
R4066 VDD.n1174 VDD.n1041 15.3605
R4067 VDD.n1184 VDD.n1041 15.3605
R4068 VDD.n1184 VDD.n1038 15.3605
R4069 VDD.n1195 VDD.n1038 15.3605
R4070 VDD.n1195 VDD.n1030 15.3605
R4071 VDD.n1206 VDD.n1030 15.3605
R4072 VDD.n1206 VDD.n1027 15.3605
R4073 VDD.n1217 VDD.n1027 15.3605
R4074 VDD.n1217 VDD.n1017 15.3605
R4075 VDD.n1231 VDD.n1017 15.3605
R4076 VDD.n1231 VDD.n1013 15.3605
R4077 VDD.n1239 VDD.n1013 15.3605
R4078 VDD.n1240 VDD.n1239 15.3605
R4079 VDD.n1241 VDD.n1240 15.3605
R4080 VDD.n800 VDD.n280 15.3605
R4081 VDD.n909 VDD.n280 15.3605
R4082 VDD.n909 VDD.n281 15.3605
R4083 VDD.n904 VDD.n281 15.3605
R4084 VDD.n904 VDD.n903 15.3605
R4085 VDD.n901 VDD.n286 15.3605
R4086 VDD.n896 VDD.n286 15.3605
R4087 VDD.n896 VDD.n895 15.3605
R4088 VDD.n895 VDD.n894 15.3605
R4089 VDD.n894 VDD.n289 15.3605
R4090 VDD.n889 VDD.n289 15.3605
R4091 VDD.n889 VDD.n888 15.3605
R4092 VDD.n888 VDD.n887 15.3605
R4093 VDD.n887 VDD.n292 15.3605
R4094 VDD.n882 VDD.n292 15.3605
R4095 VDD.n882 VDD.n881 15.3605
R4096 VDD.n881 VDD.n880 15.3605
R4097 VDD.n880 VDD.n295 15.3605
R4098 VDD.n875 VDD.n295 15.3605
R4099 VDD.n875 VDD.n874 15.3605
R4100 VDD.n874 VDD.n873 15.3605
R4101 VDD.n873 VDD.n298 15.3605
R4102 VDD.n868 VDD.n298 15.3605
R4103 VDD.n868 VDD.n867 15.3605
R4104 VDD.n867 VDD.n866 15.3605
R4105 VDD.n866 VDD.n301 15.3605
R4106 VDD.n861 VDD.n301 15.3605
R4107 VDD.n861 VDD.n860 15.3605
R4108 VDD.n860 VDD.n859 15.3605
R4109 VDD.n859 VDD.n304 15.3605
R4110 VDD.n854 VDD.n304 15.3605
R4111 VDD.n854 VDD.n853 15.3605
R4112 VDD.n853 VDD.n852 15.3605
R4113 VDD.n852 VDD.n307 15.3605
R4114 VDD.n847 VDD.n307 15.3605
R4115 VDD.n847 VDD.n846 15.3605
R4116 VDD.n846 VDD.n845 15.3605
R4117 VDD.n845 VDD.n310 15.3605
R4118 VDD.n840 VDD.n310 15.3605
R4119 VDD.n840 VDD.n839 15.3605
R4120 VDD.n839 VDD.n838 15.3605
R4121 VDD.n838 VDD.n313 15.3605
R4122 VDD.n833 VDD.n313 15.3605
R4123 VDD.n833 VDD.n832 15.3605
R4124 VDD.n832 VDD.n831 15.3605
R4125 VDD.n831 VDD.n316 15.3605
R4126 VDD.n826 VDD.n316 15.3605
R4127 VDD.n826 VDD.n825 15.3605
R4128 VDD.n825 VDD.n824 15.3605
R4129 VDD.n824 VDD.n319 15.3605
R4130 VDD.n819 VDD.n319 15.3605
R4131 VDD.n819 VDD.n818 15.3605
R4132 VDD.n818 VDD.n817 15.3605
R4133 VDD.n817 VDD.n322 15.3605
R4134 VDD.n812 VDD.n322 15.3605
R4135 VDD.n791 VDD.n325 15.3605
R4136 VDD.n810 VDD.n325 15.3605
R4137 VDD.n811 VDD.n810 15.3605
R4138 VDD.n678 VDD.n330 15.3605
R4139 VDD.n678 VDD.n677 15.3605
R4140 VDD.n684 VDD.n677 15.3605
R4141 VDD.n685 VDD.n684 15.3605
R4142 VDD.n686 VDD.n685 15.3605
R4143 VDD.n686 VDD.n675 15.3605
R4144 VDD.n692 VDD.n675 15.3605
R4145 VDD.n693 VDD.n692 15.3605
R4146 VDD.n694 VDD.n693 15.3605
R4147 VDD.n694 VDD.n673 15.3605
R4148 VDD.n700 VDD.n673 15.3605
R4149 VDD.n701 VDD.n700 15.3605
R4150 VDD.n702 VDD.n701 15.3605
R4151 VDD.n702 VDD.n671 15.3605
R4152 VDD.n708 VDD.n671 15.3605
R4153 VDD.n709 VDD.n708 15.3605
R4154 VDD.n710 VDD.n709 15.3605
R4155 VDD.n710 VDD.n669 15.3605
R4156 VDD.n716 VDD.n669 15.3605
R4157 VDD.n717 VDD.n716 15.3605
R4158 VDD.n718 VDD.n717 15.3605
R4159 VDD.n718 VDD.n667 15.3605
R4160 VDD.n724 VDD.n667 15.3605
R4161 VDD.n725 VDD.n724 15.3605
R4162 VDD.n726 VDD.n725 15.3605
R4163 VDD.n726 VDD.n665 15.3605
R4164 VDD.n732 VDD.n665 15.3605
R4165 VDD.n733 VDD.n732 15.3605
R4166 VDD.n734 VDD.n733 15.3605
R4167 VDD.n734 VDD.n663 15.3605
R4168 VDD.n740 VDD.n663 15.3605
R4169 VDD.n741 VDD.n740 15.3605
R4170 VDD.n742 VDD.n741 15.3605
R4171 VDD.n742 VDD.n661 15.3605
R4172 VDD.n748 VDD.n661 15.3605
R4173 VDD.n749 VDD.n748 15.3605
R4174 VDD.n750 VDD.n749 15.3605
R4175 VDD.n750 VDD.n659 15.3605
R4176 VDD.n756 VDD.n659 15.3605
R4177 VDD.n757 VDD.n756 15.3605
R4178 VDD.n758 VDD.n757 15.3605
R4179 VDD.n758 VDD.n657 15.3605
R4180 VDD.n764 VDD.n657 15.3605
R4181 VDD.n765 VDD.n764 15.3605
R4182 VDD.n766 VDD.n765 15.3605
R4183 VDD.n766 VDD.n655 15.3605
R4184 VDD.n772 VDD.n655 15.3605
R4185 VDD.n773 VDD.n772 15.3605
R4186 VDD.n774 VDD.n773 15.3605
R4187 VDD.n774 VDD.n653 15.3605
R4188 VDD.n780 VDD.n653 15.3605
R4189 VDD.n781 VDD.n780 15.3605
R4190 VDD.n782 VDD.n781 15.3605
R4191 VDD.n782 VDD.n651 15.3605
R4192 VDD.n651 VDD.n650 15.3605
R4193 VDD.n789 VDD.n650 15.3605
R4194 VDD.n790 VDD.n789 15.3605
R4195 VDD.n797 VDD.n796 15.3605
R4196 VDD.n806 VDD.n797 15.3605
R4197 VDD.n806 VDD.n805 15.3605
R4198 VDD.n524 VDD.n523 15.3605
R4199 VDD.n638 VDD.n524 15.3605
R4200 VDD.n638 VDD.n637 15.3605
R4201 VDD.n636 VDD.n634 15.3605
R4202 VDD.n634 VDD.n631 15.3605
R4203 VDD.n631 VDD.n630 15.3605
R4204 VDD.n630 VDD.n627 15.3605
R4205 VDD.n627 VDD.n626 15.3605
R4206 VDD.n626 VDD.n623 15.3605
R4207 VDD.n623 VDD.n622 15.3605
R4208 VDD.n622 VDD.n619 15.3605
R4209 VDD.n619 VDD.n618 15.3605
R4210 VDD.n618 VDD.n615 15.3605
R4211 VDD.n615 VDD.n614 15.3605
R4212 VDD.n614 VDD.n611 15.3605
R4213 VDD.n611 VDD.n610 15.3605
R4214 VDD.n610 VDD.n607 15.3605
R4215 VDD.n607 VDD.n606 15.3605
R4216 VDD.n606 VDD.n603 15.3605
R4217 VDD.n603 VDD.n602 15.3605
R4218 VDD.n602 VDD.n599 15.3605
R4219 VDD.n599 VDD.n598 15.3605
R4220 VDD.n598 VDD.n595 15.3605
R4221 VDD.n595 VDD.n594 15.3605
R4222 VDD.n594 VDD.n591 15.3605
R4223 VDD.n591 VDD.n590 15.3605
R4224 VDD.n590 VDD.n587 15.3605
R4225 VDD.n587 VDD.n586 15.3605
R4226 VDD.n586 VDD.n583 15.3605
R4227 VDD.n583 VDD.n582 15.3605
R4228 VDD.n582 VDD.n579 15.3605
R4229 VDD.n579 VDD.n578 15.3605
R4230 VDD.n578 VDD.n575 15.3605
R4231 VDD.n575 VDD.n574 15.3605
R4232 VDD.n574 VDD.n571 15.3605
R4233 VDD.n571 VDD.n570 15.3605
R4234 VDD.n570 VDD.n567 15.3605
R4235 VDD.n567 VDD.n566 15.3605
R4236 VDD.n566 VDD.n563 15.3605
R4237 VDD.n563 VDD.n562 15.3605
R4238 VDD.n562 VDD.n559 15.3605
R4239 VDD.n559 VDD.n558 15.3605
R4240 VDD.n558 VDD.n555 15.3605
R4241 VDD.n555 VDD.n554 15.3605
R4242 VDD.n554 VDD.n551 15.3605
R4243 VDD.n551 VDD.n550 15.3605
R4244 VDD.n550 VDD.n547 15.3605
R4245 VDD.n547 VDD.n546 15.3605
R4246 VDD.n546 VDD.n543 15.3605
R4247 VDD.n543 VDD.n542 15.3605
R4248 VDD.n542 VDD.n539 15.3605
R4249 VDD.n539 VDD.n538 15.3605
R4250 VDD.n538 VDD.n535 15.3605
R4251 VDD.n535 VDD.n534 15.3605
R4252 VDD.n534 VDD.n531 15.3605
R4253 VDD.n531 VDD.n530 15.3605
R4254 VDD.n530 VDD.n527 15.3605
R4255 VDD.n527 VDD.n526 15.3605
R4256 VDD.n526 VDD.n363 15.3605
R4257 VDD.n644 VDD.n363 15.3605
R4258 VDD.n518 VDD.n364 15.3605
R4259 VDD.n642 VDD.n364 15.3605
R4260 VDD.n643 VDD.n642 15.3605
R4261 VDD.n403 VDD.n400 15.3605
R4262 VDD.n409 VDD.n400 15.3605
R4263 VDD.n410 VDD.n409 15.3605
R4264 VDD.n413 VDD.n410 15.3605
R4265 VDD.n413 VDD.n398 15.3605
R4266 VDD.n420 VDD.n419 15.3605
R4267 VDD.n421 VDD.n420 15.3605
R4268 VDD.n421 VDD.n395 15.3605
R4269 VDD.n427 VDD.n395 15.3605
R4270 VDD.n428 VDD.n427 15.3605
R4271 VDD.n429 VDD.n428 15.3605
R4272 VDD.n429 VDD.n393 15.3605
R4273 VDD.n435 VDD.n393 15.3605
R4274 VDD.n436 VDD.n435 15.3605
R4275 VDD.n437 VDD.n436 15.3605
R4276 VDD.n437 VDD.n391 15.3605
R4277 VDD.n443 VDD.n391 15.3605
R4278 VDD.n444 VDD.n443 15.3605
R4279 VDD.n445 VDD.n444 15.3605
R4280 VDD.n445 VDD.n389 15.3605
R4281 VDD.n451 VDD.n389 15.3605
R4282 VDD.n452 VDD.n451 15.3605
R4283 VDD.n453 VDD.n452 15.3605
R4284 VDD.n453 VDD.n387 15.3605
R4285 VDD.n459 VDD.n387 15.3605
R4286 VDD.n460 VDD.n459 15.3605
R4287 VDD.n461 VDD.n460 15.3605
R4288 VDD.n461 VDD.n385 15.3605
R4289 VDD.n467 VDD.n385 15.3605
R4290 VDD.n468 VDD.n467 15.3605
R4291 VDD.n469 VDD.n468 15.3605
R4292 VDD.n469 VDD.n383 15.3605
R4293 VDD.n475 VDD.n383 15.3605
R4294 VDD.n476 VDD.n475 15.3605
R4295 VDD.n477 VDD.n476 15.3605
R4296 VDD.n477 VDD.n381 15.3605
R4297 VDD.n483 VDD.n381 15.3605
R4298 VDD.n484 VDD.n483 15.3605
R4299 VDD.n485 VDD.n484 15.3605
R4300 VDD.n485 VDD.n379 15.3605
R4301 VDD.n491 VDD.n379 15.3605
R4302 VDD.n492 VDD.n491 15.3605
R4303 VDD.n493 VDD.n492 15.3605
R4304 VDD.n493 VDD.n377 15.3605
R4305 VDD.n499 VDD.n377 15.3605
R4306 VDD.n500 VDD.n499 15.3605
R4307 VDD.n501 VDD.n500 15.3605
R4308 VDD.n501 VDD.n375 15.3605
R4309 VDD.n507 VDD.n375 15.3605
R4310 VDD.n508 VDD.n507 15.3605
R4311 VDD.n509 VDD.n508 15.3605
R4312 VDD.n509 VDD.n373 15.3605
R4313 VDD.n373 VDD.n372 15.3605
R4314 VDD.n516 VDD.n372 15.3605
R4315 VDD.n517 VDD.n516 15.3605
R4316 VDD.n207 VDD.n65 15.3605
R4317 VDD.n208 VDD.n207 15.3605
R4318 VDD.n248 VDD.n208 15.3605
R4319 VDD.n216 VDD.n215 15.3605
R4320 VDD.n222 VDD.n215 15.3605
R4321 VDD.n223 VDD.n222 15.3605
R4322 VDD.n224 VDD.n223 15.3605
R4323 VDD.n224 VDD.n213 15.3605
R4324 VDD.n230 VDD.n213 15.3605
R4325 VDD.n231 VDD.n230 15.3605
R4326 VDD.n232 VDD.n231 15.3605
R4327 VDD.n232 VDD.n211 15.3605
R4328 VDD.n238 VDD.n211 15.3605
R4329 VDD.n239 VDD.n238 15.3605
R4330 VDD.n240 VDD.n239 15.3605
R4331 VDD.n240 VDD.n209 15.3605
R4332 VDD.n246 VDD.n209 15.3605
R4333 VDD.n247 VDD.n246 15.3605
R4334 VDD.n255 VDD.n254 15.3605
R4335 VDD.n254 VDD.n253 15.3605
R4336 VDD.n253 VDD.n202 15.3605
R4337 VDD.n201 VDD.n69 15.3605
R4338 VDD.n197 VDD.n69 15.3605
R4339 VDD.n197 VDD.n196 15.3605
R4340 VDD.n196 VDD.n195 15.3605
R4341 VDD.n195 VDD.n45 15.3605
R4342 VDD.n274 VDD.n45 15.3605
R4343 VDD.n274 VDD.n273 15.3605
R4344 VDD.n273 VDD.n272 15.3605
R4345 VDD.n272 VDD.n49 15.3605
R4346 VDD.n268 VDD.n49 15.3605
R4347 VDD.n268 VDD.n267 15.3605
R4348 VDD.n267 VDD.n266 15.3605
R4349 VDD.n266 VDD.n55 15.3605
R4350 VDD.n262 VDD.n55 15.3605
R4351 VDD.n172 VDD.n83 15.3605
R4352 VDD.n121 VDD.n83 15.3605
R4353 VDD.n161 VDD.n121 15.3605
R4354 VDD.n129 VDD.n128 15.3605
R4355 VDD.n135 VDD.n128 15.3605
R4356 VDD.n136 VDD.n135 15.3605
R4357 VDD.n137 VDD.n136 15.3605
R4358 VDD.n137 VDD.n126 15.3605
R4359 VDD.n143 VDD.n126 15.3605
R4360 VDD.n144 VDD.n143 15.3605
R4361 VDD.n145 VDD.n144 15.3605
R4362 VDD.n145 VDD.n124 15.3605
R4363 VDD.n151 VDD.n124 15.3605
R4364 VDD.n152 VDD.n151 15.3605
R4365 VDD.n153 VDD.n152 15.3605
R4366 VDD.n153 VDD.n122 15.3605
R4367 VDD.n159 VDD.n122 15.3605
R4368 VDD.n160 VDD.n159 15.3605
R4369 VDD.n168 VDD.n167 15.3605
R4370 VDD.n167 VDD.n166 15.3605
R4371 VDD.n166 VDD.n116 15.3605
R4372 VDD.n112 VDD.n94 15.3605
R4373 VDD.n112 VDD.n111 15.3605
R4374 VDD.n111 VDD.n110 15.3605
R4375 VDD.n110 VDD.n108 15.3605
R4376 VDD.n108 VDD.n107 15.3605
R4377 VDD.n183 VDD.n73 15.3605
R4378 VDD.n183 VDD.n182 15.3605
R4379 VDD.n182 VDD.n181 15.3605
R4380 VDD.n181 VDD.n77 15.3605
R4381 VDD.n177 VDD.n77 15.3605
R4382 VDD.n177 VDD.n176 15.3605
R4383 VDD.n176 VDD.n175 15.3605
R4384 VDD.n521 VDD.n520 14.9939
R4385 VDD.n640 VDD.n332 14.9939
R4386 VDD.n794 VDD.n793 14.9939
R4387 VDD.n808 VDD.n327 14.9939
R4388 VDD.n1352 VDD.n920 13.2471
R4389 VDD.n1345 VDD.n1344 13.2471
R4390 VDD.n1062 VDD.n928 13.2471
R4391 VDD.n1146 VDD.n929 13.2471
R4392 VDD.n1149 VDD.n930 13.2471
R4393 VDD.n1167 VDD.n931 13.2471
R4394 VDD.n1170 VDD.n932 13.2471
R4395 VDD.n1188 VDD.n933 13.2471
R4396 VDD.n1191 VDD.n934 13.2471
R4397 VDD.n1210 VDD.n935 13.2471
R4398 VDD.n1213 VDD.n936 13.2471
R4399 VDD.n1235 VDD.n937 13.2471
R4400 VDD.n938 VDD.n937 13.2471
R4401 VDD.n1234 VDD.n936 13.2471
R4402 VDD.n1214 VDD.n935 13.2471
R4403 VDD.n1209 VDD.n934 13.2471
R4404 VDD.n1192 VDD.n933 13.2471
R4405 VDD.n1187 VDD.n932 13.2471
R4406 VDD.n1171 VDD.n931 13.2471
R4407 VDD.n1166 VDD.n930 13.2471
R4408 VDD.n1150 VDD.n929 13.2471
R4409 VDD.n1145 VDD.n928 13.2471
R4410 VDD.n1344 VDD.n927 13.2471
R4411 VDD.n926 VDD.n920 13.2471
R4412 VDD.n1353 VDD.n919 13.2471
R4413 VDD.n1397 VDD.t30 12.789
R4414 VDD.n1416 VDD.t34 12.789
R4415 VDD.n912 VDD.n911 11.8276
R4416 VDD.n1359 VDD.n913 9.40867
R4417 VDD.n1339 VDD.n941 9.40867
R4418 VDD.n1342 VDD.n1341 9.3005
R4419 VDD.n1237 VDD.n938 9.3005
R4420 VDD.n1236 VDD.n1235 9.3005
R4421 VDD.n1234 VDD.n1233 9.3005
R4422 VDD.n1213 VDD.n1016 9.3005
R4423 VDD.n1215 VDD.n1214 9.3005
R4424 VDD.n1211 VDD.n1210 9.3005
R4425 VDD.n1209 VDD.n1208 9.3005
R4426 VDD.n1191 VDD.n1029 9.3005
R4427 VDD.n1193 VDD.n1192 9.3005
R4428 VDD.n1189 VDD.n1188 9.3005
R4429 VDD.n1187 VDD.n1186 9.3005
R4430 VDD.n1170 VDD.n1040 9.3005
R4431 VDD.n1172 VDD.n1171 9.3005
R4432 VDD.n1168 VDD.n1167 9.3005
R4433 VDD.n1166 VDD.n1165 9.3005
R4434 VDD.n1149 VDD.n1051 9.3005
R4435 VDD.n1151 VDD.n1150 9.3005
R4436 VDD.n1147 VDD.n1146 9.3005
R4437 VDD.n1145 VDD.n1144 9.3005
R4438 VDD.n1063 VDD.n1062 9.3005
R4439 VDD.n1064 VDD.n927 9.3005
R4440 VDD.n1346 VDD.n1345 9.3005
R4441 VDD.n926 VDD.n921 9.3005
R4442 VDD.n1352 VDD.n1351 9.3005
R4443 VDD.n1354 VDD.n1353 9.3005
R4444 VDD.n1358 VDD.n1357 9.3005
R4445 VDD.n1356 VDD.n1355 9.3005
R4446 VDD.n918 VDD.n917 9.3005
R4447 VDD.n1350 VDD.n1349 9.3005
R4448 VDD.n1348 VDD.n1347 9.3005
R4449 VDD.n925 VDD.n924 9.3005
R4450 VDD.n1066 VDD.n1065 9.3005
R4451 VDD.n1143 VDD.n1142 9.3005
R4452 VDD.n1061 VDD.n1060 9.3005
R4453 VDD.n1153 VDD.n1152 9.3005
R4454 VDD.n1148 VDD.n1052 9.3005
R4455 VDD.n1164 VDD.n1163 9.3005
R4456 VDD.n1050 VDD.n1049 9.3005
R4457 VDD.n1174 VDD.n1173 9.3005
R4458 VDD.n1169 VDD.n1041 9.3005
R4459 VDD.n1185 VDD.n1184 9.3005
R4460 VDD.n1039 VDD.n1038 9.3005
R4461 VDD.n1195 VDD.n1194 9.3005
R4462 VDD.n1190 VDD.n1030 9.3005
R4463 VDD.n1207 VDD.n1206 9.3005
R4464 VDD.n1028 VDD.n1027 9.3005
R4465 VDD.n1217 VDD.n1216 9.3005
R4466 VDD.n1212 VDD.n1017 9.3005
R4467 VDD.n1232 VDD.n1231 9.3005
R4468 VDD.n1015 VDD.n1013 9.3005
R4469 VDD.n1239 VDD.n1238 9.3005
R4470 VDD.n1240 VDD.n939 9.3005
R4471 VDD.n280 VDD.n278 9.3005
R4472 VDD.n910 VDD.n909 9.3005
R4473 VDD.n281 VDD.n279 9.3005
R4474 VDD.n904 VDD.n285 9.3005
R4475 VDD.n411 VDD.n410 9.3005
R4476 VDD.n413 VDD.n412 9.3005
R4477 VDD.n401 VDD.n400 9.3005
R4478 VDD.n409 VDD.n277 9.3005
R4479 VDD.n270 VDD.n49 9.3005
R4480 VDD.n269 VDD.n268 9.3005
R4481 VDD.n267 VDD.n51 9.3005
R4482 VDD.n266 VDD.n265 9.3005
R4483 VDD.n264 VDD.n55 9.3005
R4484 VDD.n113 VDD.n112 9.3005
R4485 VDD.n111 VDD.n95 9.3005
R4486 VDD.n110 VDD.n109 9.3005
R4487 VDD.n108 VDD.n71 9.3005
R4488 VDD.n182 VDD.n70 9.3005
R4489 VDD.n181 VDD.n180 9.3005
R4490 VDD.n179 VDD.n77 9.3005
R4491 VDD.n178 VDD.n177 9.3005
R4492 VDD.n176 VDD.n78 9.3005
R4493 VDD.n184 VDD.n183 9.3005
R4494 VDD.n199 VDD.n69 9.3005
R4495 VDD.n198 VDD.n197 9.3005
R4496 VDD.n196 VDD.n185 9.3005
R4497 VDD.n195 VDD.n194 9.3005
R4498 VDD.n45 VDD.n42 9.3005
R4499 VDD.n201 VDD.n200 9.3005
R4500 VDD.n275 VDD.n274 9.3005
R4501 VDD.n273 VDD.n44 9.3005
R4502 VDD.n272 VDD.n271 9.3005
R4503 VDD.n1446 VDD.n17 9.3005
R4504 VDD.n1447 VDD.n1446 9.3005
R4505 VDD.n1446 VDD.n1444 9.3005
R4506 VDD.n1453 VDD.n12 9.3005
R4507 VDD.n1454 VDD.n1453 9.3005
R4508 VDD.n1453 VDD.n1452 9.3005
R4509 VDD.n1467 VDD.n1466 9.3005
R4510 VDD.n1466 VDD.n1465 9.3005
R4511 VDD.n1466 VDD.n7 9.3005
R4512 VDD.n1383 VDD.n1382 9.3005
R4513 VDD.n1366 VDD.n1363 9.3005
R4514 VDD.n1367 VDD.n1366 9.3005
R4515 VDD.n1366 VDD.n1365 9.3005
R4516 VDD.n1429 VDD.n1428 9.3005
R4517 VDD.n1429 VDD.n28 9.3005
R4518 VDD.n1430 VDD.n1429 9.3005
R4519 VDD.n1437 VDD.n27 9.3005
R4520 VDD.n1390 VDD.n1389 9.3005
R4521 VDD.n1391 VDD.n1390 9.3005
R4522 VDD.n1390 VDD.n1386 9.3005
R4523 VDD.n1427 VDD.n1426 9.3005
R4524 VDD.n1432 VDD.n1431 9.3005
R4525 VDD.n1434 VDD.n1433 9.3005
R4526 VDD.n1435 VDD.n26 9.3005
R4527 VDD.n1440 VDD.n1439 9.3005
R4528 VDD.n1441 VDD.n22 9.3005
R4529 VDD.n1443 VDD.n1442 9.3005
R4530 VDD.n21 VDD.n20 9.3005
R4531 VDD.n1449 VDD.n1448 9.3005
R4532 VDD.n1451 VDD.n1450 9.3005
R4533 VDD.n16 VDD.n15 9.3005
R4534 VDD.n1456 VDD.n1455 9.3005
R4535 VDD.n1458 VDD.n1457 9.3005
R4536 VDD.n1459 VDD.n11 9.3005
R4537 VDD.n1462 VDD.n1461 9.3005
R4538 VDD.n1464 VDD.n1463 9.3005
R4539 VDD.n8 VDD.n6 9.3005
R4540 VDD.n1468 VDD.n5 9.3005
R4541 VDD.n1470 VDD.n1469 9.3005
R4542 VDD.n1472 VDD.n1471 9.3005
R4543 VDD.n2 VDD.n0 9.3005
R4544 VDD.n1388 VDD.n32 9.3005
R4545 VDD.n1385 VDD.n36 9.3005
R4546 VDD.n1393 VDD.n1392 9.3005
R4547 VDD.n1384 VDD.n35 9.3005
R4548 VDD.n1377 VDD.n37 9.3005
R4549 VDD.n1379 VDD.n1378 9.3005
R4550 VDD.n39 VDD.n38 9.3005
R4551 VDD.n1364 VDD.n41 9.3005
R4552 VDD.n1369 VDD.n1368 9.3005
R4553 VDD.n520 VDD.t4 7.49721
R4554 VDD.n640 VDD.t4 7.49721
R4555 VDD.n793 VDD.t21 7.49721
R4556 VDD.n808 VDD.t21 7.49721
R4557 VDD.n1360 VDD.n912 6.14008
R4558 VDD.n1402 VDD.t0 5.48127
R4559 VDD.n1410 VDD.t32 5.48127
R4560 VDD.n1382 VDD.n1380 4.63585
R4561 VDD.n1438 VDD.n1437 4.63585
R4562 VDD.n1338 VDD.n943 4.26392
R4563 VDD.n1011 VDD.n940 4.26392
R4564 VDD.n263 VDD.n56 4.26392
R4565 VDD.n115 VDD.n114 4.26392
R4566 VDD.n174 VDD.n173 4.26392
R4567 VDD.n804 VDD.n798 4.25809
R4568 VDD.n902 VDD.n901 4.25809
R4569 VDD.n402 VDD.n368 4.25809
R4570 VDD.n419 VDD.n397 4.25809
R4571 VDD.n1331 VDD.n942 4.20736
R4572 VDD.n944 VDD.n942 4.20736
R4573 VDD.n107 VDD.n72 4.20736
R4574 VDD.n73 VDD.n72 4.20736
R4575 VDD.n800 VDD.n798 4.18823
R4576 VDD.n903 VDD.n902 4.18823
R4577 VDD.n398 VDD.n397 4.18823
R4578 VDD.n403 VDD.n402 4.18823
R4579 VDD.n1338 VDD.n1337 4.18603
R4580 VDD.n1241 VDD.n940 4.18603
R4581 VDD.n263 VDD.n262 4.18603
R4582 VDD.n114 VDD.n94 4.18603
R4583 VDD.n175 VDD.n174 4.18603
R4584 VDD.n200 VDD.n184 3.00131
R4585 VDD.n1343 VDD.t16 2.8655
R4586 VDD.n1363 VDD.n1362 2.78194
R4587 VDD.n264 VDD.n263 2.75514
R4588 VDD.n174 VDD.n78 2.75514
R4589 VDD.n114 VDD.n113 2.75514
R4590 VDD.n902 VDD.n285 2.73371
R4591 VDD.n798 VDD.n278 2.73371
R4592 VDD.n412 VDD.n397 2.73371
R4593 VDD.n402 VDD.n401 2.73371
R4594 VDD.n1339 VDD.n1338 2.68062
R4595 VDD.n1340 VDD.n940 2.68062
R4596 VDD.n1339 VDD.n942 2.54782
R4597 VDD.n184 VDD.n72 2.54782
R4598 VDD.n1176 VDD.t15 1.18504
R4599 VDD.n1362 VDD.n276 0.974574
R4600 VDD.n912 VDD.n277 0.410917
R4601 VDD.n1361 VDD 0.34193
R4602 VDD.n1340 VDD.n1339 0.310019
R4603 VDD.n1362 VDD.n1361 0.18325
R4604 VDD.n270 VDD.n269 0.173577
R4605 VDD.n269 VDD.n51 0.173577
R4606 VDD.n265 VDD.n51 0.173577
R4607 VDD.n265 VDD.n264 0.173577
R4608 VDD.n180 VDD.n70 0.173577
R4609 VDD.n180 VDD.n179 0.173577
R4610 VDD.n179 VDD.n178 0.173577
R4611 VDD.n178 VDD.n78 0.173577
R4612 VDD.n113 VDD.n95 0.173577
R4613 VDD.n109 VDD.n95 0.173577
R4614 VDD.n109 VDD.n71 0.173577
R4615 VDD.n184 VDD.n70 0.166365
R4616 VDD.n184 VDD.n71 0.166365
R4617 VDD.n285 VDD.n279 0.155672
R4618 VDD.n412 VDD.n411 0.155672
R4619 VDD.n910 VDD.n279 0.151025
R4620 VDD.n911 VDD.n278 0.12981
R4621 VDD.n411 VDD.n277 0.112569
R4622 VDD.n271 VDD.n270 0.105758
R4623 VDD.n1360 VDD.n1359 0.0895
R4624 VDD.n1379 VDD.n38 0.0815811
R4625 VDD.n1392 VDD.n1384 0.0815811
R4626 VDD.n1469 VDD.n1468 0.0815811
R4627 VDD.n1459 VDD.n1458 0.0815811
R4628 VDD.n1443 VDD.n22 0.0815811
R4629 VDD.n1435 VDD.n1434 0.0815811
R4630 VDD.n1389 VDD.n0 0.0739797
R4631 VDD.n1451 VDD.n17 0.0739797
R4632 VDD.n401 VDD.n277 0.0694655
R4633 VDD.n1368 VDD.n1367 0.0553986
R4634 VDD.n1383 VDD.n37 0.0553986
R4635 VDD.n1465 VDD.n1464 0.0553986
R4636 VDD.n1454 VDD.n16 0.0553986
R4637 VDD.n1439 VDD.n27 0.0553986
R4638 VDD.n1430 VDD.n1427 0.0553986
R4639 VDD.n1388 VDD.n1386 0.0537095
R4640 VDD.n1448 VDD.n1447 0.0537095
R4641 VDD.n1392 VDD.n1391 0.0486419
R4642 VDD.n1444 VDD.n1443 0.0486419
R4643 VDD.n275 VDD.n44 0.0483723
R4644 VDD.n1469 VDD.n1 0.0473536
R4645 VDD.n1460 VDD.n1459 0.0473536
R4646 VDD.n1365 VDD.n38 0.0469527
R4647 VDD.n1468 VDD.n1467 0.0469527
R4648 VDD.n1458 VDD.n12 0.0469527
R4649 VDD.n1434 VDD.n28 0.0469527
R4650 VDD.n1380 VDD.n1379 0.0456644
R4651 VDD.n1438 VDD.n1435 0.0456644
R4652 VDD.n200 VDD.n199 0.041224
R4653 VDD.n199 VDD.n198 0.041224
R4654 VDD.n198 VDD.n185 0.041224
R4655 VDD.n194 VDD.n185 0.041224
R4656 VDD.n194 VDD.n42 0.041224
R4657 VDD VDD.n0 0.0410405
R4658 VDD VDD.n1472 0.0410405
R4659 VDD.n1461 VDD 0.0410405
R4660 VDD VDD.n1451 0.0410405
R4661 VDD.n1380 VDD.n37 0.0372185
R4662 VDD.n1439 VDD.n1438 0.0372185
R4663 VDD.n1472 VDD.n1 0.0355293
R4664 VDD.n1461 VDD.n1460 0.0355293
R4665 VDD.n1365 VDD.n1364 0.0351284
R4666 VDD.n1467 VDD.n6 0.0351284
R4667 VDD VDD.n7 0.0351284
R4668 VDD.n1455 VDD.n12 0.0351284
R4669 VDD.n1452 VDD 0.0351284
R4670 VDD.n1431 VDD.n28 0.0351284
R4671 VDD.n1428 VDD 0.0351284
R4672 VDD.n1391 VDD.n1385 0.0334392
R4673 VDD.n1444 VDD.n21 0.0334392
R4674 VDD.n1386 VDD.n1385 0.0283716
R4675 VDD.n1447 VDD.n21 0.0283716
R4676 VDD.n1367 VDD.n1364 0.0266824
R4677 VDD.n1384 VDD.n1383 0.0266824
R4678 VDD.n1465 VDD.n6 0.0266824
R4679 VDD.n1455 VDD.n1454 0.0266824
R4680 VDD.n27 VDD.n22 0.0266824
R4681 VDD.n1431 VDD.n1430 0.0266824
R4682 VDD.n1361 VDD.n1360 0.026
R4683 VDD.n276 VDD.n42 0.0253869
R4684 VDD.n271 VDD.n50 0.0244362
R4685 VDD.n50 VDD.n43 0.0204468
R4686 VDD.n276 VDD.n275 0.019117
R4687 VDD.n911 VDD.n910 0.0180781
R4688 VDD.n1355 VDD.n914 0.0115063
R4689 VDD.n1354 VDD.n918 0.0115063
R4690 VDD.n1351 VDD.n1350 0.0115063
R4691 VDD.n1347 VDD.n921 0.0115063
R4692 VDD.n1346 VDD.n925 0.0115063
R4693 VDD.n1065 VDD.n1064 0.0115063
R4694 VDD.n1143 VDD.n1063 0.0115063
R4695 VDD.n1144 VDD.n1061 0.0115063
R4696 VDD.n1152 VDD.n1147 0.0115063
R4697 VDD.n1151 VDD.n1148 0.0115063
R4698 VDD.n1164 VDD.n1051 0.0115063
R4699 VDD.n1165 VDD.n1050 0.0115063
R4700 VDD.n1173 VDD.n1168 0.0115063
R4701 VDD.n1172 VDD.n1169 0.0115063
R4702 VDD.n1185 VDD.n1040 0.0115063
R4703 VDD.n1186 VDD.n1039 0.0115063
R4704 VDD.n1194 VDD.n1189 0.0115063
R4705 VDD.n1193 VDD.n1190 0.0115063
R4706 VDD.n1207 VDD.n1029 0.0115063
R4707 VDD.n1208 VDD.n1028 0.0115063
R4708 VDD.n1216 VDD.n1211 0.0115063
R4709 VDD.n1215 VDD.n1212 0.0115063
R4710 VDD.n1232 VDD.n1016 0.0115063
R4711 VDD.n1233 VDD.n1015 0.0115063
R4712 VDD.n1238 VDD.n1236 0.0115063
R4713 VDD.n1237 VDD.n939 0.0115063
R4714 VDD.n1389 VDD.n1388 0.00810135
R4715 VDD.n1448 VDD.n17 0.00810135
R4716 VDD.n276 VDD.n43 0.00790741
R4717 VDD.n1368 VDD.n1363 0.00641216
R4718 VDD.n1464 VDD.n7 0.00641216
R4719 VDD.n1452 VDD.n16 0.00641216
R4720 VDD.n1428 VDD.n1427 0.00641216
R4721 VDD.n1341 VDD.n1340 0.00505975
R4722 VDD.n1359 VDD.n1358 0.00474528
R4723 VDD.n44 VDD.n43 0.00448936
R4724 VDD.n1358 VDD.n914 0.000814465
R4725 VDD.n1355 VDD.n1354 0.000814465
R4726 VDD.n1351 VDD.n918 0.000814465
R4727 VDD.n1350 VDD.n921 0.000814465
R4728 VDD.n1347 VDD.n1346 0.000814465
R4729 VDD.n1064 VDD.n925 0.000814465
R4730 VDD.n1065 VDD.n1063 0.000814465
R4731 VDD.n1144 VDD.n1143 0.000814465
R4732 VDD.n1147 VDD.n1061 0.000814465
R4733 VDD.n1152 VDD.n1151 0.000814465
R4734 VDD.n1148 VDD.n1051 0.000814465
R4735 VDD.n1165 VDD.n1164 0.000814465
R4736 VDD.n1168 VDD.n1050 0.000814465
R4737 VDD.n1173 VDD.n1172 0.000814465
R4738 VDD.n1169 VDD.n1040 0.000814465
R4739 VDD.n1186 VDD.n1185 0.000814465
R4740 VDD.n1189 VDD.n1039 0.000814465
R4741 VDD.n1194 VDD.n1193 0.000814465
R4742 VDD.n1190 VDD.n1029 0.000814465
R4743 VDD.n1208 VDD.n1207 0.000814465
R4744 VDD.n1211 VDD.n1028 0.000814465
R4745 VDD.n1216 VDD.n1215 0.000814465
R4746 VDD.n1212 VDD.n1016 0.000814465
R4747 VDD.n1233 VDD.n1232 0.000814465
R4748 VDD.n1236 VDD.n1015 0.000814465
R4749 VDD.n1238 VDD.n1237 0.000814465
R4750 VDD.n1341 VDD.n939 0.000814465
R4751 OUT_N.n2 OUT_N.n0 272.036
R4752 OUT_N.n5 OUT_N.n3 203.779
R4753 OUT_N.n2 OUT_N.n1 181.863
R4754 OUT_N.n5 OUT_N.n4 105.144
R4755 OUT_N.n7 OUT_N.n6 29.1831
R4756 OUT_N.n4 OUT_N.t1 21.2805
R4757 OUT_N.n4 OUT_N.t0 21.2805
R4758 OUT_N.n3 OUT_N.t2 21.2805
R4759 OUT_N.n3 OUT_N.t3 21.2805
R4760 OUT_N.n1 OUT_N.t5 17.8272
R4761 OUT_N.n1 OUT_N.t4 17.8272
R4762 OUT_N.n0 OUT_N.t6 17.8272
R4763 OUT_N.n0 OUT_N.t7 17.8272
R4764 OUT_N.n6 OUT_N.n5 17.529
R4765 OUT_N.n6 OUT_N.n2 13.7643
R4766 OUT_N OUT_N.n9 12.4005
R4767 OUT_N.n9 OUT_N.n8 9.37158
R4768 OUT_N.n8 OUT_N.n7 9.36995
R4769 OUT_N.n9 OUT_N 6.8005
R4770 OUT_N.n8 OUT_N 3.27197
R4771 OUT_N OUT_N.n7 2.0005
R4772 COMP_N.n1 COMP_N.t4 448.906
R4773 COMP_N.n23 COMP_N.t3 438.723
R4774 COMP_N.n22 COMP_N.n12 285.877
R4775 COMP_N.n22 COMP_N.n13 285.877
R4776 COMP_N.n22 COMP_N.n14 285.877
R4777 COMP_N.n22 COMP_N.n15 285.877
R4778 COMP_N.n22 COMP_N.n8 292.502
R4779 COMP_N.n23 COMP_N.t5 245.976
R4780 COMP_N.n9 COMP_N.n22 14.5437
R4781 COMP_N.n17 COMP_N.n16 27.1064
R4782 COMP_N.n19 COMP_N.n18 27.1064
R4783 COMP_N.n21 COMP_N.n20 27.1064
R4784 COMP_N.n8 COMP_N.n5 29.8389
R4785 COMP_N.n8 COMP_N.n7 4.651
R4786 COMP_N.n12 COMP_N.n11 13.2471
R4787 COMP_N.n17 COMP_N.n13 13.2471
R4788 COMP_N.n19 COMP_N.n14 13.2471
R4789 COMP_N.n21 COMP_N.n15 13.2471
R4790 COMP_N.n16 COMP_N.n12 13.2471
R4791 COMP_N.n18 COMP_N.n13 13.2471
R4792 COMP_N.n20 COMP_N.n14 13.2471
R4793 COMP_N.n5 COMP_N.n15 13.2471
R4794 COMP_N.t0 COMP_N.n0 8.82296
R4795 COMP_N.n0 COMP_N.n1 0.171028
R4796 COMP_N.n6 COMP_N.n5 9.3005
R4797 COMP_N.n6 COMP_N.n21 9.3005
R4798 COMP_N.n20 COMP_N.n4 9.3005
R4799 COMP_N.n4 COMP_N.n19 9.3005
R4800 COMP_N.n18 COMP_N.n3 9.3005
R4801 COMP_N.n3 COMP_N.n17 9.3005
R4802 COMP_N.n16 COMP_N.n2 9.3005
R4803 COMP_N.n2 COMP_N.n11 9.3005
R4804 COMP_N.n9 COMP_N.n11 34.0929
R4805 COMP_N COMP_N.n10 2.48833
R4806 COMP_N.n10 COMP_N.n9 0.306732
R4807 COMP_N.n0 COMP_N.t2 18.5545
R4808 COMP_N COMP_N.n23 2.92037
R4809 COMP_N.n22 COMP_N.t1 1.433
R4810 COMP_N.n7 COMP_N.n1 0.735064
R4811 COMP_N.n10 COMP_N.n2 0.233515
R4812 COMP_N.n7 COMP_N.n6 0.231269
R4813 COMP_N.n6 COMP_N.n4 0.231269
R4814 COMP_N.n4 COMP_N.n3 0.231269
R4815 COMP_N.n3 COMP_N.n2 0.231269
R4816 a_1546_691.n1 a_1546_691.t5 448.688
R4817 a_1546_691.n51 a_1546_691.t3 438.599
R4818 a_1546_691.n95 a_1546_691.n29 285.877
R4819 a_1546_691.n95 a_1546_691.n30 285.877
R4820 a_1546_691.n95 a_1546_691.n31 285.877
R4821 a_1546_691.n95 a_1546_691.n32 285.877
R4822 a_1546_691.n95 a_1546_691.n33 285.877
R4823 a_1546_691.n95 a_1546_691.n34 285.877
R4824 a_1546_691.n95 a_1546_691.n35 285.877
R4825 a_1546_691.n95 a_1546_691.n36 285.877
R4826 a_1546_691.n95 a_1546_691.n37 285.877
R4827 a_1546_691.n95 a_1546_691.n38 285.877
R4828 a_1546_691.n95 a_1546_691.n39 285.877
R4829 a_1546_691.n95 a_1546_691.n40 285.877
R4830 a_1546_691.n95 a_1546_691.n41 285.877
R4831 a_1546_691.n95 a_1546_691.n42 285.877
R4832 a_1546_691.n95 a_1546_691.n43 285.877
R4833 a_1546_691.n95 a_1546_691.n44 285.877
R4834 a_1546_691.n95 a_1546_691.n45 285.877
R4835 a_1546_691.n95 a_1546_691.n46 285.877
R4836 a_1546_691.n95 a_1546_691.n47 285.877
R4837 a_1546_691.n95 a_1546_691.n48 285.877
R4838 a_1546_691.n95 a_1546_691.n49 285.877
R4839 a_1546_691.n95 a_1546_691.n50 285.877
R4840 a_1546_691.n95 a_1546_691.n26 292.502
R4841 a_1546_691.n51 a_1546_691.t4 246.101
R4842 a_1546_691.n1 a_1546_691.n0 0.177424
R4843 a_1546_691.n27 a_1546_691.n95 65.2288
R4844 a_1546_691.n54 a_1546_691.n53 27.1064
R4845 a_1546_691.n56 a_1546_691.n55 27.1064
R4846 a_1546_691.n58 a_1546_691.n57 27.1064
R4847 a_1546_691.n60 a_1546_691.n59 27.1064
R4848 a_1546_691.n62 a_1546_691.n61 27.1064
R4849 a_1546_691.n64 a_1546_691.n63 27.1064
R4850 a_1546_691.n66 a_1546_691.n65 27.1064
R4851 a_1546_691.n68 a_1546_691.n67 27.1064
R4852 a_1546_691.n70 a_1546_691.n69 27.1064
R4853 a_1546_691.n72 a_1546_691.n71 27.1064
R4854 a_1546_691.n74 a_1546_691.n73 27.1064
R4855 a_1546_691.n76 a_1546_691.n75 27.1064
R4856 a_1546_691.n78 a_1546_691.n77 27.1064
R4857 a_1546_691.n80 a_1546_691.n79 27.1064
R4858 a_1546_691.n82 a_1546_691.n81 27.1064
R4859 a_1546_691.n84 a_1546_691.n83 27.1064
R4860 a_1546_691.n86 a_1546_691.n85 27.1064
R4861 a_1546_691.n88 a_1546_691.n87 27.1064
R4862 a_1546_691.n90 a_1546_691.n89 27.1064
R4863 a_1546_691.n92 a_1546_691.n91 27.1064
R4864 a_1546_691.n94 a_1546_691.n93 27.1064
R4865 a_1546_691.n26 a_1546_691.n23 29.8389
R4866 a_1546_691.n26 a_1546_691.n25 4.651
R4867 a_1546_691.n52 a_1546_691.n29 13.2471
R4868 a_1546_691.n54 a_1546_691.n30 13.2471
R4869 a_1546_691.n56 a_1546_691.n31 13.2471
R4870 a_1546_691.n58 a_1546_691.n32 13.2471
R4871 a_1546_691.n60 a_1546_691.n33 13.2471
R4872 a_1546_691.n62 a_1546_691.n34 13.2471
R4873 a_1546_691.n64 a_1546_691.n35 13.2471
R4874 a_1546_691.n66 a_1546_691.n36 13.2471
R4875 a_1546_691.n68 a_1546_691.n37 13.2471
R4876 a_1546_691.n70 a_1546_691.n38 13.2471
R4877 a_1546_691.n72 a_1546_691.n39 13.2471
R4878 a_1546_691.n74 a_1546_691.n40 13.2471
R4879 a_1546_691.n76 a_1546_691.n41 13.2471
R4880 a_1546_691.n78 a_1546_691.n42 13.2471
R4881 a_1546_691.n80 a_1546_691.n43 13.2471
R4882 a_1546_691.n82 a_1546_691.n44 13.2471
R4883 a_1546_691.n84 a_1546_691.n45 13.2471
R4884 a_1546_691.n86 a_1546_691.n46 13.2471
R4885 a_1546_691.n88 a_1546_691.n47 13.2471
R4886 a_1546_691.n90 a_1546_691.n48 13.2471
R4887 a_1546_691.n92 a_1546_691.n49 13.2471
R4888 a_1546_691.n94 a_1546_691.n50 13.2471
R4889 a_1546_691.n53 a_1546_691.n29 13.2471
R4890 a_1546_691.n55 a_1546_691.n30 13.2471
R4891 a_1546_691.n57 a_1546_691.n31 13.2471
R4892 a_1546_691.n59 a_1546_691.n32 13.2471
R4893 a_1546_691.n61 a_1546_691.n33 13.2471
R4894 a_1546_691.n63 a_1546_691.n34 13.2471
R4895 a_1546_691.n65 a_1546_691.n35 13.2471
R4896 a_1546_691.n67 a_1546_691.n36 13.2471
R4897 a_1546_691.n69 a_1546_691.n37 13.2471
R4898 a_1546_691.n71 a_1546_691.n38 13.2471
R4899 a_1546_691.n73 a_1546_691.n39 13.2471
R4900 a_1546_691.n75 a_1546_691.n40 13.2471
R4901 a_1546_691.n77 a_1546_691.n41 13.2471
R4902 a_1546_691.n79 a_1546_691.n42 13.2471
R4903 a_1546_691.n81 a_1546_691.n43 13.2471
R4904 a_1546_691.n83 a_1546_691.n44 13.2471
R4905 a_1546_691.n85 a_1546_691.n45 13.2471
R4906 a_1546_691.n87 a_1546_691.n46 13.2471
R4907 a_1546_691.n89 a_1546_691.n47 13.2471
R4908 a_1546_691.n91 a_1546_691.n48 13.2471
R4909 a_1546_691.n93 a_1546_691.n49 13.2471
R4910 a_1546_691.n23 a_1546_691.n50 13.2471
R4911 a_1546_691.n1 a_1546_691.t0 18.3315
R4912 a_1546_691.n24 a_1546_691.n23 9.3005
R4913 a_1546_691.n24 a_1546_691.n94 9.3005
R4914 a_1546_691.n93 a_1546_691.n22 9.3005
R4915 a_1546_691.n22 a_1546_691.n92 9.3005
R4916 a_1546_691.n91 a_1546_691.n21 9.3005
R4917 a_1546_691.n21 a_1546_691.n90 9.3005
R4918 a_1546_691.n89 a_1546_691.n20 9.3005
R4919 a_1546_691.n20 a_1546_691.n88 9.3005
R4920 a_1546_691.n87 a_1546_691.n19 9.3005
R4921 a_1546_691.n19 a_1546_691.n86 9.3005
R4922 a_1546_691.n85 a_1546_691.n18 9.3005
R4923 a_1546_691.n18 a_1546_691.n84 9.3005
R4924 a_1546_691.n83 a_1546_691.n17 9.3005
R4925 a_1546_691.n17 a_1546_691.n82 9.3005
R4926 a_1546_691.n81 a_1546_691.n16 9.3005
R4927 a_1546_691.n16 a_1546_691.n80 9.3005
R4928 a_1546_691.n79 a_1546_691.n15 9.3005
R4929 a_1546_691.n15 a_1546_691.n78 9.3005
R4930 a_1546_691.n77 a_1546_691.n14 9.3005
R4931 a_1546_691.n14 a_1546_691.n76 9.3005
R4932 a_1546_691.n75 a_1546_691.n13 9.3005
R4933 a_1546_691.n13 a_1546_691.n74 9.3005
R4934 a_1546_691.n73 a_1546_691.n12 9.3005
R4935 a_1546_691.n12 a_1546_691.n72 9.3005
R4936 a_1546_691.n71 a_1546_691.n11 9.3005
R4937 a_1546_691.n11 a_1546_691.n70 9.3005
R4938 a_1546_691.n69 a_1546_691.n10 9.3005
R4939 a_1546_691.n10 a_1546_691.n68 9.3005
R4940 a_1546_691.n67 a_1546_691.n9 9.3005
R4941 a_1546_691.n9 a_1546_691.n66 9.3005
R4942 a_1546_691.n65 a_1546_691.n8 9.3005
R4943 a_1546_691.n8 a_1546_691.n64 9.3005
R4944 a_1546_691.n63 a_1546_691.n7 9.3005
R4945 a_1546_691.n7 a_1546_691.n62 9.3005
R4946 a_1546_691.n61 a_1546_691.n6 9.3005
R4947 a_1546_691.n6 a_1546_691.n60 9.3005
R4948 a_1546_691.n59 a_1546_691.n5 9.3005
R4949 a_1546_691.n5 a_1546_691.n58 9.3005
R4950 a_1546_691.n57 a_1546_691.n4 9.3005
R4951 a_1546_691.n4 a_1546_691.n56 9.3005
R4952 a_1546_691.n55 a_1546_691.n3 9.3005
R4953 a_1546_691.n3 a_1546_691.n54 9.3005
R4954 a_1546_691.n53 a_1546_691.n2 9.3005
R4955 a_1546_691.n2 a_1546_691.n52 9.3005
R4956 a_1546_691.n52 a_1546_691.n27 33.3013
R4957 a_1546_691.n51 a_1546_691.n28 6.1339
R4958 a_1546_691.n27 a_1546_691.n28 1.11007
R4959 a_1546_691.n0 a_1546_691.t1 8.81146
R4960 a_1546_691.t2 a_1546_691.n95 1.433
R4961 a_1546_691.n25 a_1546_691.n0 0.99182
R4962 a_1546_691.n25 a_1546_691.n24 0.231269
R4963 a_1546_691.n24 a_1546_691.n22 0.231269
R4964 a_1546_691.n22 a_1546_691.n21 0.231269
R4965 a_1546_691.n21 a_1546_691.n20 0.231269
R4966 a_1546_691.n20 a_1546_691.n19 0.231269
R4967 a_1546_691.n19 a_1546_691.n18 0.231269
R4968 a_1546_691.n18 a_1546_691.n17 0.231269
R4969 a_1546_691.n17 a_1546_691.n16 0.231269
R4970 a_1546_691.n16 a_1546_691.n15 0.231269
R4971 a_1546_691.n15 a_1546_691.n14 0.231269
R4972 a_1546_691.n14 a_1546_691.n13 0.231269
R4973 a_1546_691.n13 a_1546_691.n12 0.231269
R4974 a_1546_691.n12 a_1546_691.n11 0.231269
R4975 a_1546_691.n11 a_1546_691.n10 0.231269
R4976 a_1546_691.n10 a_1546_691.n9 0.231269
R4977 a_1546_691.n9 a_1546_691.n8 0.231269
R4978 a_1546_691.n8 a_1546_691.n7 0.231269
R4979 a_1546_691.n7 a_1546_691.n6 0.231269
R4980 a_1546_691.n6 a_1546_691.n5 0.231269
R4981 a_1546_691.n5 a_1546_691.n4 0.231269
R4982 a_1546_691.n4 a_1546_691.n3 0.231269
R4983 a_1546_691.n3 a_1546_691.n2 0.231269
R4984 a_1546_691.n28 a_1546_691.n2 0.230249
R4985 IN_P IN_P.t0 1166.07
R4986 CLK CLK.t0 683.186
R4987 IN_N IN_N.t0 1164.84
C0 VDD IN_N 0.492526f
C1 VDD SR_set 1.71377f
C2 sky130_fd_sc_hvl__nand2_1_0.A sky130_fd_sc_hvl__buf_4$VAR1_0.A 0.42053f
C3 sky130_fd_sc_hvl__nand2_1_0.A SR_reset 0.268426f
C4 sky130_fd_sc_hvl__buf_4$VAR1_0.A OUT_N 0.017328f
C5 IN_P COMP_N 0.505271f
C6 sky130_fd_sc_hvl__nand2_1_0.A OUT_P 0.022293f
C7 VDD a_6094_6197# 0.948432f
C8 VDD a_6094_4183# 0.961465f
C9 sky130_fd_sc_hvl__buf_4$VAR1_0.A SR_reset 0.101739f
C10 OUT_P SR_reset 0.012198f
C11 sky130_fd_sc_hvl__nand2_1_0.A SR_set 0.106395f
C12 SR_set OUT_N 0.023572f
C13 IN_N IN_P 0.3836f
C14 sky130_fd_sc_hvl__nand2_1_0.A a_6094_6197# 0.353494f
C15 SR_set COMP_N 0.508972f
C16 VDD CLK 0.056711f
C17 a_6094_4183# OUT_N 0.643433f
C18 SR_set sky130_fd_sc_hvl__buf_4$VAR1_0.A 0.174424f
C19 SR_set SR_reset 0.070561f
C20 a_6094_4183# sky130_fd_sc_hvl__buf_4$VAR1_0.A 0.265631f
C21 SR_reset a_6094_6197# 0.060205f
C22 OUT_P a_6094_6197# 0.643767f
C23 VDD sky130_fd_sc_hvl__nand2_1_0.A 0.93545f
C24 VDD OUT_N 0.830496f
C25 VDD COMP_N 2.46865f
C26 VDD IN_P 0.576344f
C27 CLK COMP_N 0.426329f
C28 VDD sky130_fd_sc_hvl__buf_4$VAR1_0.A 0.957821f
C29 SR_set a_6094_4183# 0.052234f
C30 VDD SR_reset 1.87486f
C31 VDD OUT_P 0.83212f
C32 CLK VSS 1.23452f
C33 OUT_N VSS 1.09356f
C34 OUT_P VSS 1.10172f
C35 IN_P VSS 0.63687f
C36 IN_N VSS 0.532662f
C37 VDD VSS 63.93357f
C38 a_6094_4183# VSS 1.43951f
C39 SR_set VSS 2.29631f
C40 sky130_fd_sc_hvl__buf_4$VAR1_0.A VSS 1.01393f
C41 sky130_fd_sc_hvl__nand2_1_0.A VSS 0.918837f
C42 a_6094_6197# VSS 1.37358f
C43 SR_reset VSS 2.00343f
C44 COMP_N VSS 6.092555f
C45 a_1546_691.n0 VSS 1.13556f
C46 a_1546_691.n1 VSS 1.93353f
C47 a_1546_691.n2 VSS 0.034159f
C48 a_1546_691.n3 VSS 0.032611f
C49 a_1546_691.n4 VSS 0.032611f
C50 a_1546_691.n5 VSS 0.032611f
C51 a_1546_691.n6 VSS 0.032611f
C52 a_1546_691.n7 VSS 0.032611f
C53 a_1546_691.n8 VSS 0.032611f
C54 a_1546_691.n9 VSS 0.032611f
C55 a_1546_691.n10 VSS 0.032611f
C56 a_1546_691.n11 VSS 0.032611f
C57 a_1546_691.n12 VSS 0.032611f
C58 a_1546_691.n13 VSS 0.032611f
C59 a_1546_691.n14 VSS 0.032611f
C60 a_1546_691.n15 VSS 0.032611f
C61 a_1546_691.n16 VSS 0.032611f
C62 a_1546_691.n17 VSS 0.032611f
C63 a_1546_691.n18 VSS 0.032611f
C64 a_1546_691.n19 VSS 0.032611f
C65 a_1546_691.n20 VSS 0.032611f
C66 a_1546_691.n21 VSS 0.032611f
C67 a_1546_691.n22 VSS 0.032611f
C68 a_1546_691.n24 VSS 0.032611f
C69 a_1546_691.n25 VSS 0.483077f
C70 a_1546_691.n27 VSS 0.022194f
C71 a_1546_691.n28 VSS 0.450893f
C72 a_1546_691.t1 VSS 0.30663f
C73 a_1546_691.t0 VSS 0.153403f
C74 a_1546_691.t5 VSS 0.254486f
C75 a_1546_691.t4 VSS 0.065992f
C76 a_1546_691.t3 VSS 0.251331f
C77 a_1546_691.n51 VSS 0.501274f
C78 a_1546_691.n95 VSS 0.524225f
C79 a_1546_691.t2 VSS 0.174206f
C80 COMP_N.n0 VSS 0.853184f
C81 COMP_N.n1 VSS 1.48497f
C82 COMP_N.n2 VSS 0.023604f
C83 COMP_N.n3 VSS 0.022154f
C84 COMP_N.n4 VSS 0.022154f
C85 COMP_N.n6 VSS 0.022154f
C86 COMP_N.n7 VSS 0.071249f
C87 COMP_N.n9 VSS 0.159464f
C88 COMP_N.n10 VSS 0.497555f
C89 COMP_N.t0 VSS 0.210161f
C90 COMP_N.t2 VSS 0.115282f
C91 COMP_N.t4 VSS 0.17305f
C92 COMP_N.t1 VSS 0.118346f
C93 COMP_N.n22 VSS 0.433115f
C94 COMP_N.t5 VSS 0.044801f
C95 COMP_N.t3 VSS 0.170765f
C96 COMP_N.n23 VSS 0.191281f
C97 VDD.n1 VSS 0.024158f
C98 VDD.t36 VSS 0.013666f
C99 VDD.t30 VSS 0.013666f
C100 VDD.n33 VSS 0.016086f
C101 VDD.t7 VSS 0.033246f
C102 VDD.t18 VSS 0.03048f
C103 VDD.n50 VSS 0.054515f
C104 VDD.n63 VSS 0.156935f
C105 VDD.n66 VSS 0.046182f
C106 VDD.t3 VSS 0.030564f
C107 VDD.n90 VSS 0.156935f
C108 VDD.n91 VSS 0.046182f
C109 VDD.t2 VSS 0.030788f
C110 VDD.n119 VSS 0.156935f
C111 VDD.n163 VSS 0.08253f
C112 VDD.n164 VSS 0.046182f
C113 VDD.n170 VSS 0.08253f
C114 VDD.n184 VSS 0.213165f
C115 VDD.n200 VSS 0.164807f
C116 VDD.t17 VSS 0.030788f
C117 VDD.n205 VSS 0.156935f
C118 VDD.n250 VSS 0.08253f
C119 VDD.n251 VSS 0.046182f
C120 VDD.n257 VSS 0.08253f
C121 VDD.n276 VSS 0.160804f
C122 VDD.n283 VSS 0.458346f
C123 VDD.t21 VSS 0.089921f
C124 VDD.n327 VSS 0.241037f
C125 VDD.n332 VSS 0.241037f
C126 VDD.t4 VSS 0.089921f
C127 VDD.n370 VSS 0.458346f
C128 VDD.n520 VSS 0.134881f
C129 VDD.n521 VSS 0.241037f
C130 VDD.n640 VSS 0.134881f
C131 VDD.n647 VSS 0.458346f
C132 VDD.n648 VSS 0.458346f
C133 VDD.n793 VSS 0.134881f
C134 VDD.n794 VSS 0.241037f
C135 VDD.n808 VSS 0.134881f
C136 VDD.n911 VSS 0.024809f
C137 VDD.n912 VSS 0.076256f
C138 VDD.n914 VSS 0.016425f
C139 VDD.n918 VSS 0.01567f
C140 VDD.n921 VSS 0.01567f
C141 VDD.n925 VSS 0.01567f
C142 VDD.t16 VSS 0.016426f
C143 VDD.n939 VSS 0.01567f
C144 VDD.n947 VSS 0.081675f
C145 VDD.n951 VSS 0.081675f
C146 VDD.n965 VSS 0.081675f
C147 VDD.n979 VSS 0.063232f
C148 VDD.n1015 VSS 0.01567f
C149 VDD.n1016 VSS 0.01567f
C150 VDD.n1020 VSS 0.063232f
C151 VDD.n1025 VSS 0.063232f
C152 VDD.n1028 VSS 0.01567f
C153 VDD.n1029 VSS 0.01567f
C154 VDD.n1032 VSS 0.063232f
C155 VDD.n1036 VSS 0.063232f
C156 VDD.n1039 VSS 0.01567f
C157 VDD.n1040 VSS 0.01567f
C158 VDD.n1043 VSS 0.062354f
C159 VDD.n1047 VSS 0.063232f
C160 VDD.t15 VSS 0.031616f
C161 VDD.n1050 VSS 0.01567f
C162 VDD.n1051 VSS 0.01567f
C163 VDD.n1054 VSS 0.063232f
C164 VDD.n1058 VSS 0.063232f
C165 VDD.n1061 VSS 0.01567f
C166 VDD.n1063 VSS 0.01567f
C167 VDD.n1064 VSS 0.01567f
C168 VDD.n1065 VSS 0.01567f
C169 VDD.n1068 VSS 0.063232f
C170 VDD.n1073 VSS 0.063232f
C171 VDD.n1077 VSS 0.158081f
C172 VDD.n1123 VSS 0.081675f
C173 VDD.n1124 VSS 0.063232f
C174 VDD.n1125 VSS 0.063232f
C175 VDD.n1131 VSS 0.063232f
C176 VDD.n1132 VSS 0.063232f
C177 VDD.n1134 VSS 0.063232f
C178 VDD.n1140 VSS 0.063232f
C179 VDD.n1143 VSS 0.01567f
C180 VDD.n1144 VSS 0.01567f
C181 VDD.n1147 VSS 0.01567f
C182 VDD.n1148 VSS 0.01567f
C183 VDD.n1151 VSS 0.01567f
C184 VDD.n1152 VSS 0.01567f
C185 VDD.n1155 VSS 0.063232f
C186 VDD.n1161 VSS 0.063232f
C187 VDD.n1164 VSS 0.01567f
C188 VDD.n1165 VSS 0.01567f
C189 VDD.n1168 VSS 0.01567f
C190 VDD.n1169 VSS 0.01567f
C191 VDD.n1172 VSS 0.01567f
C192 VDD.n1173 VSS 0.01567f
C193 VDD.n1176 VSS 0.032494f
C194 VDD.n1182 VSS 0.063232f
C195 VDD.n1185 VSS 0.01567f
C196 VDD.n1186 VSS 0.01567f
C197 VDD.n1189 VSS 0.01567f
C198 VDD.n1190 VSS 0.01567f
C199 VDD.n1193 VSS 0.01567f
C200 VDD.n1194 VSS 0.01567f
C201 VDD.n1197 VSS 0.063232f
C202 VDD.n1204 VSS 0.063232f
C203 VDD.n1207 VSS 0.01567f
C204 VDD.n1208 VSS 0.01567f
C205 VDD.n1211 VSS 0.01567f
C206 VDD.n1212 VSS 0.01567f
C207 VDD.n1215 VSS 0.01567f
C208 VDD.n1216 VSS 0.01567f
C209 VDD.n1219 VSS 0.063232f
C210 VDD.n1227 VSS 0.063232f
C211 VDD.n1228 VSS 0.063232f
C212 VDD.n1229 VSS 0.063232f
C213 VDD.n1232 VSS 0.01567f
C214 VDD.n1233 VSS 0.01567f
C215 VDD.n1236 VSS 0.01567f
C216 VDD.n1237 VSS 0.01567f
C217 VDD.n1238 VSS 0.01567f
C218 VDD.n1243 VSS 0.063232f
C219 VDD.n1249 VSS 0.158081f
C220 VDD.n1288 VSS 0.158081f
C221 VDD.n1328 VSS 0.158081f
C222 VDD.n1333 VSS 0.048302f
C223 VDD.t13 VSS 0.031616f
C224 VDD.n1334 VSS 0.046546f
C225 VDD.n1335 VSS 0.063232f
C226 VDD.n1339 VSS 0.152209f
C227 VDD.n1340 VSS 0.192945f
C228 VDD.n1343 VSS 0.049277f
C229 VDD.n1346 VSS 0.01567f
C230 VDD.n1347 VSS 0.01567f
C231 VDD.n1350 VSS 0.01567f
C232 VDD.n1351 VSS 0.01567f
C233 VDD.n1354 VSS 0.01567f
C234 VDD.n1355 VSS 0.01567f
C235 VDD.n1359 VSS 0.056752f
C236 VDD.n1360 VSS 0.111278f
C237 VDD.n1361 VSS 3.38217f
C238 VDD.n1362 VSS 1.02162f
C239 VDD.n1363 VSS 0.214315f
C240 VDD.n1366 VSS 0.035414f
C241 VDD.n1369 VSS 0.011956f
C242 VDD.n1370 VSS 0.039657f
C243 VDD.n1373 VSS 0.019503f
C244 VDD.n1374 VSS 0.016371f
C245 VDD.t11 VSS 0.013666f
C246 VDD.t9 VSS 0.013666f
C247 VDD.n1375 VSS 0.022208f
C248 VDD.n1382 VSS 0.030238f
C249 VDD.n1390 VSS 0.029366f
C250 VDD.n1395 VSS 0.019787f
C251 VDD.t5 VSS 0.013666f
C252 VDD.n1396 VSS 0.021211f
C253 VDD.n1397 VSS 0.014663f
C254 VDD.n1400 VSS 0.026336f
C255 VDD.n1401 VSS 0.026905f
C256 VDD.t0 VSS 0.013666f
C257 VDD.n1402 VSS 0.014093f
C258 VDD.n1403 VSS 0.02178f
C259 VDD.n1406 VSS 0.019218f
C260 VDD.n1407 VSS 0.027332f
C261 VDD.n1408 VSS 0.026905f
C262 VDD.t32 VSS 0.013666f
C263 VDD.n1410 VSS 0.014093f
C264 VDD.n1411 VSS 0.02178f
C265 VDD.t19 VSS 0.013666f
C266 VDD.n1412 VSS 0.019218f
C267 VDD.n1414 VSS 0.027332f
C268 VDD.n1415 VSS 0.026336f
C269 VDD.t34 VSS 0.013666f
C270 VDD.n1416 VSS 0.014663f
C271 VDD.n1418 VSS 0.021211f
C272 VDD.t26 VSS 0.013666f
C273 VDD.n1419 VSS 0.019787f
C274 VDD.n1420 VSS 0.016086f
C275 VDD.t28 VSS 0.013666f
C276 VDD.n1421 VSS 0.022208f
C277 VDD.t24 VSS 0.013666f
C278 VDD.n1423 VSS 0.016371f
C279 VDD.n1424 VSS 0.019503f
C280 VDD.t22 VSS 0.033246f
C281 VDD.n1425 VSS 0.039657f
C282 VDD.n1426 VSS 0.011956f
C283 VDD.n1429 VSS 0.035414f
C284 VDD.n1437 VSS 0.030238f
C285 VDD.n1446 VSS 0.029366f
C286 VDD.n1453 VSS 0.035414f
C287 VDD.n1460 VSS 0.024158f
C288 VDD.n1466 VSS 0.035414f
C289 a_1077_8251.n0 VSS 1.4985f
C290 a_1077_8251.n1 VSS 1.85272f
C291 a_1077_8251.n4 VSS 1.85272f
C292 a_1077_8251.n7 VSS 3.19957f
C293 a_1077_8251.n36 VSS 0.492732f
C294 a_1077_8251.t1 VSS 0.315915f
C295 a_1077_8251.t2 VSS 0.163552f
C296 a_1077_8251.n73 VSS 0.492732f
C297 a_1077_8251.t0 VSS 0.163552f
C298 a_84_7283.n0 VSS 0.063478f
C299 a_84_7283.n3 VSS 0.012696f
C300 a_84_7283.n5 VSS 0.063478f
C301 a_84_7283.n7 VSS 0.012696f
C302 a_84_7283.n9 VSS 0.063478f
C303 a_84_7283.t0 VSS 0.182981f
C304 a_84_7283.n11 VSS 0.089521f
C305 a_84_7283.n13 VSS 0.063478f
C306 a_84_7283.t3 VSS 2.42866f
C307 a_84_7283.n15 VSS 0.012696f
C308 a_84_7283.n17 VSS 0.063478f
C309 a_84_7283.n19 VSS 0.028537f
C310 a_84_7283.n21 VSS 0.063478f
C311 a_84_7283.n23 VSS 0.0645f
C312 a_84_7283.n26 VSS 0.063478f
C313 a_84_7283.n29 VSS 0.028537f
C314 a_84_7283.n30 VSS 0.012696f
C315 a_84_7283.n32 VSS 0.063478f
C316 a_84_7283.n34 VSS 0.012696f
C317 a_84_7283.n35 VSS 0.012696f
C318 a_84_7283.n37 VSS 0.012696f
C319 a_84_7283.n39 VSS 0.063478f
C320 a_84_7283.n41 VSS 0.012696f
C321 a_84_7283.n43 VSS 0.838081f
C322 a_84_7283.n46 VSS 0.063478f
C323 a_84_7283.n49 VSS 0.012696f
C324 a_84_7283.n50 VSS 0.012696f
C325 a_84_7283.n52 VSS 0.063478f
C326 a_84_7283.n54 VSS 0.012696f
C327 a_84_7283.n55 VSS 0.012696f
C328 a_84_7283.n56 VSS 0.028537f
C329 a_84_7283.n59 VSS 0.063478f
C330 a_84_7283.n61 VSS 0.028537f
C331 a_84_7283.n63 VSS 0.110019f
C332 a_84_7283.t1 VSS 0.01743f
C333 a_84_7283.n64 VSS 0.282224f
C334 a_84_7283.t2 VSS 0.785931f
.ends

